// This is the unpowered netlist.
module caravel_hack_soc (wb_clk_i,
    wb_rst_i,
    wbs_ack_o,
    wbs_cyc_i,
    wbs_stb_i,
    wbs_we_i,
    io_in,
    io_oeb,
    io_out,
    irq,
    la_data_in,
    la_data_out,
    la_oenb,
    wbs_adr_i,
    wbs_dat_i,
    wbs_dat_o,
    wbs_sel_i);
 input wb_clk_i;
 input wb_rst_i;
 output wbs_ack_o;
 input wbs_cyc_i;
 input wbs_stb_i;
 input wbs_we_i;
 input [37:0] io_in;
 output [37:0] io_oeb;
 output [37:0] io_out;
 output [2:0] irq;
 input [63:0] la_data_in;
 output [63:0] la_data_out;
 input [63:0] la_oenb;
 input [31:0] wbs_adr_i;
 input [31:0] wbs_dat_i;
 output [31:0] wbs_dat_o;
 input [3:0] wbs_sel_i;

 wire _00000_;
 wire _00001_;
 wire _00002_;
 wire _00003_;
 wire _00004_;
 wire _00005_;
 wire _00006_;
 wire _00007_;
 wire _00008_;
 wire _00009_;
 wire _00010_;
 wire _00011_;
 wire _00012_;
 wire _00013_;
 wire _00014_;
 wire _00015_;
 wire _00016_;
 wire _00017_;
 wire _00018_;
 wire _00019_;
 wire _00020_;
 wire _00021_;
 wire _00022_;
 wire _00023_;
 wire _00024_;
 wire _00025_;
 wire _00026_;
 wire _00027_;
 wire _00028_;
 wire _00029_;
 wire _00030_;
 wire _00031_;
 wire _00032_;
 wire _00033_;
 wire _00034_;
 wire _00035_;
 wire _00036_;
 wire _00037_;
 wire _00038_;
 wire _00039_;
 wire _00040_;
 wire _00041_;
 wire _00042_;
 wire _00043_;
 wire _00044_;
 wire _00045_;
 wire _00046_;
 wire _00047_;
 wire _00048_;
 wire _00049_;
 wire _00050_;
 wire _00051_;
 wire _00052_;
 wire _00053_;
 wire _00054_;
 wire _00055_;
 wire _00056_;
 wire _00057_;
 wire _00058_;
 wire _00059_;
 wire _00060_;
 wire _00061_;
 wire _00062_;
 wire _00063_;
 wire _00064_;
 wire _00065_;
 wire _00066_;
 wire _00067_;
 wire _00068_;
 wire _00069_;
 wire _00070_;
 wire _00071_;
 wire _00072_;
 wire _00073_;
 wire _00074_;
 wire _00075_;
 wire _00076_;
 wire _00077_;
 wire _00078_;
 wire _00079_;
 wire _00080_;
 wire _00081_;
 wire _00082_;
 wire _00083_;
 wire _00084_;
 wire _00085_;
 wire _00086_;
 wire _00087_;
 wire _00088_;
 wire _00089_;
 wire _00090_;
 wire _00091_;
 wire _00092_;
 wire _00093_;
 wire _00094_;
 wire _00095_;
 wire _00096_;
 wire _00097_;
 wire _00098_;
 wire _00099_;
 wire _00100_;
 wire _00101_;
 wire _00102_;
 wire _00103_;
 wire _00104_;
 wire _00105_;
 wire _00106_;
 wire _00107_;
 wire _00108_;
 wire _00109_;
 wire _00110_;
 wire _00111_;
 wire _00112_;
 wire _00113_;
 wire _00114_;
 wire _00115_;
 wire _00116_;
 wire _00117_;
 wire _00118_;
 wire _00119_;
 wire _00120_;
 wire _00121_;
 wire _00122_;
 wire _00123_;
 wire _00124_;
 wire _00125_;
 wire _00126_;
 wire _00127_;
 wire _00128_;
 wire _00129_;
 wire _00130_;
 wire _00131_;
 wire _00132_;
 wire _00133_;
 wire _00134_;
 wire _00135_;
 wire _00136_;
 wire _00137_;
 wire _00138_;
 wire _00139_;
 wire _00140_;
 wire _00141_;
 wire _00142_;
 wire _00143_;
 wire _00144_;
 wire _00145_;
 wire _00146_;
 wire _00147_;
 wire _00148_;
 wire _00149_;
 wire _00150_;
 wire _00151_;
 wire _00152_;
 wire _00153_;
 wire _00154_;
 wire _00155_;
 wire _00156_;
 wire _00157_;
 wire _00158_;
 wire _00159_;
 wire _00160_;
 wire _00161_;
 wire _00162_;
 wire _00163_;
 wire _00164_;
 wire _00165_;
 wire _00166_;
 wire _00167_;
 wire _00168_;
 wire _00169_;
 wire _00170_;
 wire _00171_;
 wire _00172_;
 wire _00173_;
 wire _00174_;
 wire _00175_;
 wire _00176_;
 wire _00177_;
 wire _00178_;
 wire _00179_;
 wire _00180_;
 wire _00181_;
 wire _00182_;
 wire _00183_;
 wire _00184_;
 wire _00185_;
 wire _00186_;
 wire _00187_;
 wire _00188_;
 wire _00189_;
 wire _00190_;
 wire _00191_;
 wire _00192_;
 wire _00193_;
 wire _00194_;
 wire _00195_;
 wire _00196_;
 wire _00197_;
 wire _00198_;
 wire _00199_;
 wire _00200_;
 wire _00201_;
 wire _00202_;
 wire _00203_;
 wire _00204_;
 wire _00205_;
 wire _00206_;
 wire _00207_;
 wire _00208_;
 wire _00209_;
 wire _00210_;
 wire _00211_;
 wire _00212_;
 wire _00213_;
 wire _00214_;
 wire _00215_;
 wire _00216_;
 wire _00217_;
 wire _00218_;
 wire _00219_;
 wire _00220_;
 wire _00221_;
 wire _00222_;
 wire _00223_;
 wire _00224_;
 wire _00225_;
 wire _00226_;
 wire _00227_;
 wire _00228_;
 wire _00229_;
 wire _00230_;
 wire _00231_;
 wire _00232_;
 wire _00233_;
 wire _00234_;
 wire _00235_;
 wire _00236_;
 wire _00237_;
 wire _00238_;
 wire _00239_;
 wire _00240_;
 wire _00241_;
 wire _00242_;
 wire _00243_;
 wire _00244_;
 wire _00245_;
 wire _00246_;
 wire _00247_;
 wire _00248_;
 wire _00249_;
 wire _00250_;
 wire _00251_;
 wire _00252_;
 wire _00253_;
 wire _00254_;
 wire _00255_;
 wire _00256_;
 wire _00257_;
 wire _00258_;
 wire _00259_;
 wire _00260_;
 wire _00261_;
 wire _00262_;
 wire _00263_;
 wire _00264_;
 wire _00265_;
 wire _00266_;
 wire _00267_;
 wire _00268_;
 wire _00269_;
 wire _00270_;
 wire _00271_;
 wire _00272_;
 wire _00273_;
 wire _00274_;
 wire _00275_;
 wire _00276_;
 wire _00277_;
 wire _00278_;
 wire _00279_;
 wire _00280_;
 wire _00281_;
 wire _00282_;
 wire _00283_;
 wire _00284_;
 wire _00285_;
 wire _00286_;
 wire _00287_;
 wire _00288_;
 wire _00289_;
 wire _00290_;
 wire _00291_;
 wire _00292_;
 wire _00293_;
 wire _00294_;
 wire _00295_;
 wire _00296_;
 wire _00297_;
 wire _00298_;
 wire _00299_;
 wire _00300_;
 wire _00301_;
 wire _00302_;
 wire _00303_;
 wire _00304_;
 wire _00305_;
 wire _00306_;
 wire _00307_;
 wire _00308_;
 wire _00309_;
 wire _00310_;
 wire _00311_;
 wire _00312_;
 wire _00313_;
 wire _00314_;
 wire _00315_;
 wire _00316_;
 wire _00317_;
 wire _00318_;
 wire _00319_;
 wire _00320_;
 wire _00321_;
 wire _00322_;
 wire _00323_;
 wire _00324_;
 wire _00325_;
 wire _00326_;
 wire _00327_;
 wire _00328_;
 wire _00329_;
 wire _00330_;
 wire _00331_;
 wire _00332_;
 wire _00333_;
 wire _00334_;
 wire _00335_;
 wire _00336_;
 wire _00337_;
 wire _00338_;
 wire _00339_;
 wire _00340_;
 wire _00341_;
 wire _00342_;
 wire _00343_;
 wire _00344_;
 wire _00345_;
 wire _00346_;
 wire _00347_;
 wire _00348_;
 wire _00349_;
 wire _00350_;
 wire _00351_;
 wire _00352_;
 wire _00353_;
 wire _00354_;
 wire _00355_;
 wire _00356_;
 wire _00357_;
 wire _00358_;
 wire _00359_;
 wire _00360_;
 wire _00361_;
 wire _00362_;
 wire _00363_;
 wire _00364_;
 wire _00365_;
 wire _00366_;
 wire _00367_;
 wire _00368_;
 wire _00369_;
 wire _00370_;
 wire _00371_;
 wire _00372_;
 wire _00373_;
 wire _00374_;
 wire _00375_;
 wire _00376_;
 wire _00377_;
 wire _00378_;
 wire _00379_;
 wire _00380_;
 wire _00381_;
 wire _00382_;
 wire _00383_;
 wire _00384_;
 wire _00385_;
 wire _00386_;
 wire _00387_;
 wire _00388_;
 wire _00389_;
 wire _00390_;
 wire _00391_;
 wire _00392_;
 wire _00393_;
 wire _00394_;
 wire _00395_;
 wire _00396_;
 wire _00397_;
 wire _00398_;
 wire _00399_;
 wire _00400_;
 wire _00401_;
 wire _00402_;
 wire _00403_;
 wire _00404_;
 wire _00405_;
 wire _00406_;
 wire _00407_;
 wire _00408_;
 wire _00409_;
 wire _00410_;
 wire _00411_;
 wire _00412_;
 wire _00413_;
 wire _00414_;
 wire _00415_;
 wire _00416_;
 wire _00417_;
 wire _00418_;
 wire _00419_;
 wire _00420_;
 wire _00421_;
 wire _00422_;
 wire _00423_;
 wire _00424_;
 wire _00425_;
 wire _00426_;
 wire _00427_;
 wire _00428_;
 wire _00429_;
 wire _00430_;
 wire _00431_;
 wire _00432_;
 wire _00433_;
 wire _00434_;
 wire _00435_;
 wire _00436_;
 wire _00437_;
 wire _00438_;
 wire _00439_;
 wire _00440_;
 wire _00441_;
 wire _00442_;
 wire _00443_;
 wire _00444_;
 wire _00445_;
 wire _00446_;
 wire _00447_;
 wire _00448_;
 wire _00449_;
 wire _00450_;
 wire _00451_;
 wire _00452_;
 wire _00453_;
 wire _00454_;
 wire _00455_;
 wire _00456_;
 wire _00457_;
 wire _00458_;
 wire _00459_;
 wire _00460_;
 wire _00461_;
 wire _00462_;
 wire _00463_;
 wire _00464_;
 wire _00465_;
 wire _00466_;
 wire _00467_;
 wire _00468_;
 wire _00469_;
 wire _00470_;
 wire _00471_;
 wire _00472_;
 wire _00473_;
 wire _00474_;
 wire _00475_;
 wire _00476_;
 wire _00477_;
 wire _00478_;
 wire _00479_;
 wire _00480_;
 wire _00481_;
 wire _00482_;
 wire _00483_;
 wire _00484_;
 wire _00485_;
 wire _00486_;
 wire _00487_;
 wire _00488_;
 wire _00489_;
 wire _00490_;
 wire _00491_;
 wire _00492_;
 wire _00493_;
 wire _00494_;
 wire _00495_;
 wire _00496_;
 wire _00497_;
 wire _00498_;
 wire _00499_;
 wire _00500_;
 wire _00501_;
 wire _00502_;
 wire _00503_;
 wire _00504_;
 wire _00505_;
 wire _00506_;
 wire _00507_;
 wire _00508_;
 wire _00509_;
 wire _00510_;
 wire _00511_;
 wire _00512_;
 wire _00513_;
 wire _00514_;
 wire _00515_;
 wire _00516_;
 wire _00517_;
 wire _00518_;
 wire _00519_;
 wire _00520_;
 wire _00521_;
 wire _00522_;
 wire _00523_;
 wire _00524_;
 wire _00525_;
 wire _00526_;
 wire _00527_;
 wire _00528_;
 wire _00529_;
 wire _00530_;
 wire _00531_;
 wire _00532_;
 wire _00533_;
 wire _00534_;
 wire _00535_;
 wire _00536_;
 wire _00537_;
 wire _00538_;
 wire _00539_;
 wire _00540_;
 wire _00541_;
 wire _00542_;
 wire _00543_;
 wire _00544_;
 wire _00545_;
 wire _00546_;
 wire _00547_;
 wire _00548_;
 wire _00549_;
 wire _00550_;
 wire _00551_;
 wire _00552_;
 wire _00553_;
 wire _00554_;
 wire _00555_;
 wire _00556_;
 wire _00557_;
 wire _00558_;
 wire _00559_;
 wire _00560_;
 wire _00561_;
 wire _00562_;
 wire _00563_;
 wire _00564_;
 wire _00565_;
 wire _00566_;
 wire _00567_;
 wire _00568_;
 wire _00569_;
 wire _00570_;
 wire _00571_;
 wire _00572_;
 wire _00573_;
 wire _00574_;
 wire _00575_;
 wire _00576_;
 wire _00577_;
 wire _00578_;
 wire _00579_;
 wire _00580_;
 wire _00581_;
 wire _00582_;
 wire _00583_;
 wire _00584_;
 wire _00585_;
 wire _00586_;
 wire _00587_;
 wire _00588_;
 wire _00589_;
 wire _00590_;
 wire _00591_;
 wire _00592_;
 wire _00593_;
 wire _00594_;
 wire _00595_;
 wire _00596_;
 wire _00597_;
 wire _00598_;
 wire _00599_;
 wire _00600_;
 wire _00601_;
 wire _00602_;
 wire _00603_;
 wire _00604_;
 wire _00605_;
 wire _00606_;
 wire _00607_;
 wire _00608_;
 wire _00609_;
 wire _00610_;
 wire _00611_;
 wire _00612_;
 wire _00613_;
 wire _00614_;
 wire _00615_;
 wire _00616_;
 wire _00617_;
 wire _00618_;
 wire _00619_;
 wire _00620_;
 wire _00621_;
 wire _00622_;
 wire _00623_;
 wire _00624_;
 wire _00625_;
 wire _00626_;
 wire _00627_;
 wire _00628_;
 wire _00629_;
 wire _00630_;
 wire _00631_;
 wire _00632_;
 wire _00633_;
 wire _00634_;
 wire _00635_;
 wire _00636_;
 wire _00637_;
 wire _00638_;
 wire _00639_;
 wire _00640_;
 wire _00641_;
 wire _00642_;
 wire _00643_;
 wire _00644_;
 wire _00645_;
 wire _00646_;
 wire _00647_;
 wire _00648_;
 wire _00649_;
 wire _00650_;
 wire _00651_;
 wire _00652_;
 wire _00653_;
 wire _00654_;
 wire _00655_;
 wire _00656_;
 wire _00657_;
 wire _00658_;
 wire _00659_;
 wire _00660_;
 wire _00661_;
 wire _00662_;
 wire _00663_;
 wire _00664_;
 wire _00665_;
 wire _00666_;
 wire _00667_;
 wire _00668_;
 wire _00669_;
 wire _00670_;
 wire _00671_;
 wire _00672_;
 wire _00673_;
 wire _00674_;
 wire _00675_;
 wire _00676_;
 wire _00677_;
 wire _00678_;
 wire _00679_;
 wire _00680_;
 wire _00681_;
 wire _00682_;
 wire _00683_;
 wire _00684_;
 wire _00685_;
 wire _00686_;
 wire _00687_;
 wire _00688_;
 wire _00689_;
 wire _00690_;
 wire _00691_;
 wire _00692_;
 wire _00693_;
 wire _00694_;
 wire _00695_;
 wire _00696_;
 wire _00697_;
 wire _00698_;
 wire _00699_;
 wire _00700_;
 wire _00701_;
 wire _00702_;
 wire _00703_;
 wire _00704_;
 wire _00705_;
 wire _00706_;
 wire _00707_;
 wire _00708_;
 wire _00709_;
 wire _00710_;
 wire _00711_;
 wire _00712_;
 wire _00713_;
 wire _00714_;
 wire _00715_;
 wire _00716_;
 wire _00717_;
 wire _00718_;
 wire _00719_;
 wire _00720_;
 wire _00721_;
 wire _00722_;
 wire _00723_;
 wire _00724_;
 wire _00725_;
 wire _00726_;
 wire _00727_;
 wire _00728_;
 wire _00729_;
 wire _00730_;
 wire _00731_;
 wire _00732_;
 wire _00733_;
 wire _00734_;
 wire _00735_;
 wire _00736_;
 wire _00737_;
 wire _00738_;
 wire _00739_;
 wire _00740_;
 wire _00741_;
 wire _00742_;
 wire _00743_;
 wire _00744_;
 wire _00745_;
 wire _00746_;
 wire _00747_;
 wire _00748_;
 wire _00749_;
 wire _00750_;
 wire _00751_;
 wire _00752_;
 wire _00753_;
 wire _00754_;
 wire _00755_;
 wire _00756_;
 wire _00757_;
 wire _00758_;
 wire _00759_;
 wire _00760_;
 wire _00761_;
 wire _00762_;
 wire _00763_;
 wire _00764_;
 wire _00765_;
 wire _00766_;
 wire _00767_;
 wire _00768_;
 wire _00769_;
 wire _00770_;
 wire _00771_;
 wire _00772_;
 wire _00773_;
 wire _00774_;
 wire _00775_;
 wire _00776_;
 wire _00777_;
 wire _00778_;
 wire _00779_;
 wire _00780_;
 wire _00781_;
 wire _00782_;
 wire _00783_;
 wire _00784_;
 wire _00785_;
 wire _00786_;
 wire _00787_;
 wire _00788_;
 wire _00789_;
 wire _00790_;
 wire _00791_;
 wire _00792_;
 wire _00793_;
 wire _00794_;
 wire _00795_;
 wire _00796_;
 wire _00797_;
 wire _00798_;
 wire _00799_;
 wire _00800_;
 wire _00801_;
 wire _00802_;
 wire _00803_;
 wire _00804_;
 wire _00805_;
 wire _00806_;
 wire _00807_;
 wire _00808_;
 wire _00809_;
 wire _00810_;
 wire _00811_;
 wire _00812_;
 wire _00813_;
 wire _00814_;
 wire _00815_;
 wire _00816_;
 wire _00817_;
 wire _00818_;
 wire _00819_;
 wire _00820_;
 wire _00821_;
 wire _00822_;
 wire _00823_;
 wire _00824_;
 wire _00825_;
 wire _00826_;
 wire _00827_;
 wire _00828_;
 wire _00829_;
 wire _00830_;
 wire _00831_;
 wire _00832_;
 wire _00833_;
 wire _00834_;
 wire _00835_;
 wire _00836_;
 wire _00837_;
 wire _00838_;
 wire _00839_;
 wire _00840_;
 wire _00841_;
 wire _00842_;
 wire _00843_;
 wire _00844_;
 wire _00845_;
 wire _00846_;
 wire _00847_;
 wire _00848_;
 wire _00849_;
 wire _00850_;
 wire _00851_;
 wire _00852_;
 wire _00853_;
 wire _00854_;
 wire _00855_;
 wire _00856_;
 wire _00857_;
 wire _00858_;
 wire _00859_;
 wire _00860_;
 wire _00861_;
 wire _00862_;
 wire _00863_;
 wire _00864_;
 wire _00865_;
 wire _00866_;
 wire _00867_;
 wire _00868_;
 wire _00869_;
 wire _00870_;
 wire _00871_;
 wire _00872_;
 wire _00873_;
 wire _00874_;
 wire _00875_;
 wire _00876_;
 wire _00877_;
 wire _00878_;
 wire _00879_;
 wire _00880_;
 wire _00881_;
 wire _00882_;
 wire _00883_;
 wire _00884_;
 wire _00885_;
 wire _00886_;
 wire _00887_;
 wire _00888_;
 wire _00889_;
 wire _00890_;
 wire _00891_;
 wire _00892_;
 wire _00893_;
 wire _00894_;
 wire _00895_;
 wire _00896_;
 wire _00897_;
 wire _00898_;
 wire _00899_;
 wire _00900_;
 wire _00901_;
 wire _00902_;
 wire _00903_;
 wire _00904_;
 wire _00905_;
 wire _00906_;
 wire _00907_;
 wire _00908_;
 wire _00909_;
 wire _00910_;
 wire _00911_;
 wire _00912_;
 wire _00913_;
 wire _00914_;
 wire _00915_;
 wire _00916_;
 wire _00917_;
 wire _00918_;
 wire _00919_;
 wire _00920_;
 wire _00921_;
 wire _00922_;
 wire _00923_;
 wire _00924_;
 wire _00925_;
 wire _00926_;
 wire _00927_;
 wire _00928_;
 wire _00929_;
 wire _00930_;
 wire _00931_;
 wire _00932_;
 wire _00933_;
 wire _00934_;
 wire _00935_;
 wire _00936_;
 wire _00937_;
 wire _00938_;
 wire _00939_;
 wire _00940_;
 wire _00941_;
 wire _00942_;
 wire _00943_;
 wire _00944_;
 wire _00945_;
 wire _00946_;
 wire _00947_;
 wire _00948_;
 wire _00949_;
 wire _00950_;
 wire _00951_;
 wire _00952_;
 wire _00953_;
 wire _00954_;
 wire _00955_;
 wire _00956_;
 wire _00957_;
 wire _00958_;
 wire _00959_;
 wire _00960_;
 wire _00961_;
 wire _00962_;
 wire _00963_;
 wire _00964_;
 wire _00965_;
 wire _00966_;
 wire _00967_;
 wire _00968_;
 wire _00969_;
 wire _00970_;
 wire _00971_;
 wire _00972_;
 wire _00973_;
 wire _00974_;
 wire _00975_;
 wire _00976_;
 wire _00977_;
 wire _00978_;
 wire _00979_;
 wire _00980_;
 wire _00981_;
 wire _00982_;
 wire _00983_;
 wire _00984_;
 wire _00985_;
 wire _00986_;
 wire _00987_;
 wire _00988_;
 wire _00989_;
 wire _00990_;
 wire _00991_;
 wire _00992_;
 wire _00993_;
 wire _00994_;
 wire _00995_;
 wire _00996_;
 wire _00997_;
 wire _00998_;
 wire _00999_;
 wire _01000_;
 wire _01001_;
 wire _01002_;
 wire _01003_;
 wire _01004_;
 wire _01005_;
 wire _01006_;
 wire _01007_;
 wire _01008_;
 wire _01009_;
 wire _01010_;
 wire _01011_;
 wire _01012_;
 wire _01013_;
 wire _01014_;
 wire _01015_;
 wire _01016_;
 wire _01017_;
 wire _01018_;
 wire _01019_;
 wire _01020_;
 wire _01021_;
 wire _01022_;
 wire _01023_;
 wire _01024_;
 wire _01025_;
 wire _01026_;
 wire _01027_;
 wire _01028_;
 wire _01029_;
 wire _01030_;
 wire _01031_;
 wire _01032_;
 wire _01033_;
 wire _01034_;
 wire _01035_;
 wire _01036_;
 wire _01037_;
 wire _01038_;
 wire _01039_;
 wire _01040_;
 wire _01041_;
 wire _01042_;
 wire _01043_;
 wire _01044_;
 wire _01045_;
 wire _01046_;
 wire _01047_;
 wire _01048_;
 wire _01049_;
 wire _01050_;
 wire _01051_;
 wire _01052_;
 wire _01053_;
 wire _01054_;
 wire _01055_;
 wire _01056_;
 wire _01057_;
 wire _01058_;
 wire _01059_;
 wire _01060_;
 wire _01061_;
 wire _01062_;
 wire _01063_;
 wire _01064_;
 wire _01065_;
 wire _01066_;
 wire _01067_;
 wire _01068_;
 wire _01069_;
 wire _01070_;
 wire _01071_;
 wire _01072_;
 wire _01073_;
 wire _01074_;
 wire _01075_;
 wire _01076_;
 wire _01077_;
 wire _01078_;
 wire _01079_;
 wire _01080_;
 wire _01081_;
 wire _01082_;
 wire _01083_;
 wire _01084_;
 wire _01085_;
 wire _01086_;
 wire _01087_;
 wire _01088_;
 wire _01089_;
 wire _01090_;
 wire _01091_;
 wire _01092_;
 wire _01093_;
 wire _01094_;
 wire _01095_;
 wire _01096_;
 wire _01097_;
 wire _01098_;
 wire _01099_;
 wire _01100_;
 wire _01101_;
 wire _01102_;
 wire _01103_;
 wire _01104_;
 wire _01105_;
 wire _01106_;
 wire _01107_;
 wire _01108_;
 wire _01109_;
 wire _01110_;
 wire _01111_;
 wire _01112_;
 wire _01113_;
 wire _01114_;
 wire _01115_;
 wire _01116_;
 wire _01117_;
 wire _01118_;
 wire _01119_;
 wire _01120_;
 wire _01121_;
 wire _01122_;
 wire _01123_;
 wire _01124_;
 wire _01125_;
 wire _01126_;
 wire _01127_;
 wire _01128_;
 wire _01129_;
 wire _01130_;
 wire _01131_;
 wire _01132_;
 wire _01133_;
 wire _01134_;
 wire _01135_;
 wire _01136_;
 wire _01137_;
 wire _01138_;
 wire _01139_;
 wire _01140_;
 wire _01141_;
 wire _01142_;
 wire _01143_;
 wire _01144_;
 wire _01145_;
 wire _01146_;
 wire _01147_;
 wire _01148_;
 wire _01149_;
 wire _01150_;
 wire _01151_;
 wire _01152_;
 wire _01153_;
 wire _01154_;
 wire _01155_;
 wire _01156_;
 wire _01157_;
 wire _01158_;
 wire _01159_;
 wire _01160_;
 wire _01161_;
 wire _01162_;
 wire _01163_;
 wire _01164_;
 wire _01165_;
 wire _01166_;
 wire _01167_;
 wire _01168_;
 wire _01169_;
 wire _01170_;
 wire _01171_;
 wire _01172_;
 wire _01173_;
 wire _01174_;
 wire _01175_;
 wire _01176_;
 wire _01177_;
 wire _01178_;
 wire _01179_;
 wire _01180_;
 wire _01181_;
 wire _01182_;
 wire _01183_;
 wire _01184_;
 wire _01185_;
 wire _01186_;
 wire _01187_;
 wire _01188_;
 wire _01189_;
 wire _01190_;
 wire _01191_;
 wire _01192_;
 wire _01193_;
 wire _01194_;
 wire _01195_;
 wire _01196_;
 wire _01197_;
 wire _01198_;
 wire _01199_;
 wire _01200_;
 wire _01201_;
 wire _01202_;
 wire _01203_;
 wire _01204_;
 wire _01205_;
 wire _01206_;
 wire _01207_;
 wire _01208_;
 wire _01209_;
 wire _01210_;
 wire _01211_;
 wire _01212_;
 wire _01213_;
 wire _01214_;
 wire _01215_;
 wire _01216_;
 wire _01217_;
 wire _01218_;
 wire _01219_;
 wire _01220_;
 wire _01221_;
 wire _01222_;
 wire _01223_;
 wire _01224_;
 wire _01225_;
 wire _01226_;
 wire _01227_;
 wire _01228_;
 wire _01229_;
 wire _01230_;
 wire _01231_;
 wire _01232_;
 wire _01233_;
 wire _01234_;
 wire _01235_;
 wire _01236_;
 wire _01237_;
 wire _01238_;
 wire _01239_;
 wire _01240_;
 wire _01241_;
 wire _01242_;
 wire _01243_;
 wire _01244_;
 wire _01245_;
 wire _01246_;
 wire _01247_;
 wire _01248_;
 wire _01249_;
 wire _01250_;
 wire _01251_;
 wire _01252_;
 wire _01253_;
 wire _01254_;
 wire _01255_;
 wire _01256_;
 wire _01257_;
 wire _01258_;
 wire _01259_;
 wire _01260_;
 wire _01261_;
 wire _01262_;
 wire _01263_;
 wire _01264_;
 wire _01265_;
 wire _01266_;
 wire _01267_;
 wire _01268_;
 wire _01269_;
 wire _01270_;
 wire _01271_;
 wire _01272_;
 wire _01273_;
 wire _01274_;
 wire _01275_;
 wire _01276_;
 wire _01277_;
 wire _01278_;
 wire _01279_;
 wire _01280_;
 wire _01281_;
 wire _01282_;
 wire _01283_;
 wire _01284_;
 wire _01285_;
 wire _01286_;
 wire _01287_;
 wire _01288_;
 wire _01289_;
 wire _01290_;
 wire _01291_;
 wire _01292_;
 wire _01293_;
 wire _01294_;
 wire _01295_;
 wire _01296_;
 wire _01297_;
 wire _01298_;
 wire _01299_;
 wire _01300_;
 wire _01301_;
 wire _01302_;
 wire _01303_;
 wire _01304_;
 wire _01305_;
 wire _01306_;
 wire _01307_;
 wire _01308_;
 wire _01309_;
 wire _01310_;
 wire _01311_;
 wire _01312_;
 wire _01313_;
 wire _01314_;
 wire _01315_;
 wire _01316_;
 wire _01317_;
 wire _01318_;
 wire _01319_;
 wire _01320_;
 wire _01321_;
 wire _01322_;
 wire _01323_;
 wire _01324_;
 wire _01325_;
 wire _01326_;
 wire _01327_;
 wire _01328_;
 wire _01329_;
 wire _01330_;
 wire _01331_;
 wire _01332_;
 wire _01333_;
 wire _01334_;
 wire _01335_;
 wire _01336_;
 wire _01337_;
 wire _01338_;
 wire _01339_;
 wire _01340_;
 wire _01341_;
 wire _01342_;
 wire _01343_;
 wire _01344_;
 wire _01345_;
 wire _01346_;
 wire _01347_;
 wire _01348_;
 wire _01349_;
 wire _01350_;
 wire _01351_;
 wire _01352_;
 wire _01353_;
 wire _01354_;
 wire _01355_;
 wire _01356_;
 wire _01357_;
 wire _01358_;
 wire _01359_;
 wire _01360_;
 wire _01361_;
 wire _01362_;
 wire _01363_;
 wire _01364_;
 wire _01365_;
 wire _01366_;
 wire _01367_;
 wire _01368_;
 wire _01369_;
 wire _01370_;
 wire _01371_;
 wire _01372_;
 wire _01373_;
 wire _01374_;
 wire _01375_;
 wire _01376_;
 wire _01377_;
 wire _01378_;
 wire _01379_;
 wire _01380_;
 wire _01381_;
 wire _01382_;
 wire _01383_;
 wire _01384_;
 wire _01385_;
 wire _01386_;
 wire _01387_;
 wire _01388_;
 wire _01389_;
 wire _01390_;
 wire _01391_;
 wire _01392_;
 wire _01393_;
 wire _01394_;
 wire _01395_;
 wire _01396_;
 wire _01397_;
 wire _01398_;
 wire _01399_;
 wire _01400_;
 wire _01401_;
 wire _01402_;
 wire _01403_;
 wire _01404_;
 wire _01405_;
 wire _01406_;
 wire _01407_;
 wire _01408_;
 wire _01409_;
 wire _01410_;
 wire _01411_;
 wire _01412_;
 wire _01413_;
 wire _01414_;
 wire _01415_;
 wire _01416_;
 wire _01417_;
 wire _01418_;
 wire _01419_;
 wire _01420_;
 wire _01421_;
 wire _01422_;
 wire _01423_;
 wire _01424_;
 wire _01425_;
 wire _01426_;
 wire _01427_;
 wire _01428_;
 wire _01429_;
 wire _01430_;
 wire _01431_;
 wire _01432_;
 wire _01433_;
 wire _01434_;
 wire _01435_;
 wire _01436_;
 wire _01437_;
 wire _01438_;
 wire _01439_;
 wire _01440_;
 wire _01441_;
 wire _01442_;
 wire _01443_;
 wire _01444_;
 wire _01445_;
 wire _01446_;
 wire _01447_;
 wire _01448_;
 wire _01449_;
 wire _01450_;
 wire _01451_;
 wire _01452_;
 wire _01453_;
 wire _01454_;
 wire _01455_;
 wire _01456_;
 wire _01457_;
 wire _01458_;
 wire _01459_;
 wire _01460_;
 wire _01461_;
 wire _01462_;
 wire _01463_;
 wire _01464_;
 wire _01465_;
 wire _01466_;
 wire _01467_;
 wire _01468_;
 wire _01469_;
 wire _01470_;
 wire _01471_;
 wire _01472_;
 wire _01473_;
 wire _01474_;
 wire _01475_;
 wire _01476_;
 wire _01477_;
 wire _01478_;
 wire _01479_;
 wire _01480_;
 wire _01481_;
 wire _01482_;
 wire _01483_;
 wire _01484_;
 wire _01485_;
 wire _01486_;
 wire _01487_;
 wire _01488_;
 wire _01489_;
 wire _01490_;
 wire _01491_;
 wire _01492_;
 wire _01493_;
 wire _01494_;
 wire _01495_;
 wire _01496_;
 wire _01497_;
 wire _01498_;
 wire _01499_;
 wire _01500_;
 wire _01501_;
 wire _01502_;
 wire _01503_;
 wire _01504_;
 wire _01505_;
 wire _01506_;
 wire _01507_;
 wire _01508_;
 wire _01509_;
 wire _01510_;
 wire _01511_;
 wire _01512_;
 wire _01513_;
 wire _01514_;
 wire _01515_;
 wire _01516_;
 wire _01517_;
 wire _01518_;
 wire _01519_;
 wire _01520_;
 wire _01521_;
 wire _01522_;
 wire _01523_;
 wire _01524_;
 wire _01525_;
 wire _01526_;
 wire _01527_;
 wire _01528_;
 wire _01529_;
 wire _01530_;
 wire _01531_;
 wire _01532_;
 wire _01533_;
 wire _01534_;
 wire _01535_;
 wire _01536_;
 wire _01537_;
 wire _01538_;
 wire _01539_;
 wire _01540_;
 wire _01541_;
 wire _01542_;
 wire _01543_;
 wire _01544_;
 wire _01545_;
 wire _01546_;
 wire _01547_;
 wire _01548_;
 wire _01549_;
 wire _01550_;
 wire _01551_;
 wire _01552_;
 wire _01553_;
 wire _01554_;
 wire _01555_;
 wire _01556_;
 wire _01557_;
 wire _01558_;
 wire _01559_;
 wire _01560_;
 wire _01561_;
 wire _01562_;
 wire _01563_;
 wire _01564_;
 wire _01565_;
 wire _01566_;
 wire _01567_;
 wire _01568_;
 wire _01569_;
 wire _01570_;
 wire _01571_;
 wire _01572_;
 wire _01573_;
 wire _01574_;
 wire _01575_;
 wire _01576_;
 wire _01577_;
 wire _01578_;
 wire _01579_;
 wire _01580_;
 wire _01581_;
 wire _01582_;
 wire _01583_;
 wire _01584_;
 wire _01585_;
 wire _01586_;
 wire _01587_;
 wire _01588_;
 wire _01589_;
 wire _01590_;
 wire _01591_;
 wire _01592_;
 wire _01593_;
 wire _01594_;
 wire _01595_;
 wire _01596_;
 wire _01597_;
 wire _01598_;
 wire _01599_;
 wire _01600_;
 wire _01601_;
 wire _01602_;
 wire _01603_;
 wire _01604_;
 wire _01605_;
 wire _01606_;
 wire _01607_;
 wire _01608_;
 wire _01609_;
 wire _01610_;
 wire _01611_;
 wire _01612_;
 wire _01613_;
 wire _01614_;
 wire _01615_;
 wire _01616_;
 wire _01617_;
 wire _01618_;
 wire _01619_;
 wire _01620_;
 wire _01621_;
 wire _01622_;
 wire _01623_;
 wire _01624_;
 wire _01625_;
 wire _01626_;
 wire _01627_;
 wire _01628_;
 wire _01629_;
 wire _01630_;
 wire _01631_;
 wire _01632_;
 wire _01633_;
 wire _01634_;
 wire _01635_;
 wire _01636_;
 wire _01637_;
 wire _01638_;
 wire _01639_;
 wire _01640_;
 wire _01641_;
 wire _01642_;
 wire _01643_;
 wire _01644_;
 wire _01645_;
 wire _01646_;
 wire _01647_;
 wire _01648_;
 wire _01649_;
 wire _01650_;
 wire _01651_;
 wire _01652_;
 wire _01653_;
 wire _01654_;
 wire _01655_;
 wire _01656_;
 wire _01657_;
 wire _01658_;
 wire _01659_;
 wire _01660_;
 wire _01661_;
 wire _01662_;
 wire _01663_;
 wire _01664_;
 wire _01665_;
 wire _01666_;
 wire _01667_;
 wire _01668_;
 wire _01669_;
 wire _01670_;
 wire _01671_;
 wire _01672_;
 wire _01673_;
 wire _01674_;
 wire _01675_;
 wire _01676_;
 wire _01677_;
 wire _01678_;
 wire _01679_;
 wire _01680_;
 wire _01681_;
 wire _01682_;
 wire _01683_;
 wire _01684_;
 wire _01685_;
 wire _01686_;
 wire _01687_;
 wire _01688_;
 wire _01689_;
 wire _01690_;
 wire _01691_;
 wire _01692_;
 wire _01693_;
 wire _01694_;
 wire _01695_;
 wire _01696_;
 wire _01697_;
 wire _01698_;
 wire _01699_;
 wire _01700_;
 wire _01701_;
 wire _01702_;
 wire _01703_;
 wire _01704_;
 wire _01705_;
 wire _01706_;
 wire _01707_;
 wire _01708_;
 wire _01709_;
 wire _01710_;
 wire _01711_;
 wire _01712_;
 wire _01713_;
 wire _01714_;
 wire _01715_;
 wire _01716_;
 wire _01717_;
 wire _01718_;
 wire _01719_;
 wire _01720_;
 wire _01721_;
 wire _01722_;
 wire _01723_;
 wire _01724_;
 wire _01725_;
 wire _01726_;
 wire _01727_;
 wire _01728_;
 wire _01729_;
 wire _01730_;
 wire _01731_;
 wire _01732_;
 wire _01733_;
 wire _01734_;
 wire _01735_;
 wire _01736_;
 wire _01737_;
 wire _01738_;
 wire _01739_;
 wire _01740_;
 wire _01741_;
 wire _01742_;
 wire _01743_;
 wire _01744_;
 wire _01745_;
 wire _01746_;
 wire _01747_;
 wire _01748_;
 wire _01749_;
 wire _01750_;
 wire _01751_;
 wire _01752_;
 wire _01753_;
 wire _01754_;
 wire _01755_;
 wire _01756_;
 wire _01757_;
 wire _01758_;
 wire _01759_;
 wire _01760_;
 wire _01761_;
 wire _01762_;
 wire _01763_;
 wire _01764_;
 wire _01765_;
 wire _01766_;
 wire _01767_;
 wire _01768_;
 wire _01769_;
 wire _01770_;
 wire _01771_;
 wire _01772_;
 wire _01773_;
 wire _01774_;
 wire _01775_;
 wire _01776_;
 wire _01777_;
 wire _01778_;
 wire _01779_;
 wire _01780_;
 wire _01781_;
 wire _01782_;
 wire _01783_;
 wire _01784_;
 wire _01785_;
 wire _01786_;
 wire _01787_;
 wire _01788_;
 wire _01789_;
 wire _01790_;
 wire _01791_;
 wire _01792_;
 wire _01793_;
 wire _01794_;
 wire _01795_;
 wire _01796_;
 wire _01797_;
 wire _01798_;
 wire _01799_;
 wire _01800_;
 wire _01801_;
 wire _01802_;
 wire _01803_;
 wire _01804_;
 wire _01805_;
 wire _01806_;
 wire _01807_;
 wire _01808_;
 wire _01809_;
 wire _01810_;
 wire _01811_;
 wire _01812_;
 wire _01813_;
 wire _01814_;
 wire _01815_;
 wire _01816_;
 wire _01817_;
 wire _01818_;
 wire _01819_;
 wire _01820_;
 wire _01821_;
 wire _01822_;
 wire _01823_;
 wire _01824_;
 wire _01825_;
 wire _01826_;
 wire _01827_;
 wire _01828_;
 wire _01829_;
 wire _01830_;
 wire _01831_;
 wire _01832_;
 wire _01833_;
 wire _01834_;
 wire _01835_;
 wire _01836_;
 wire _01837_;
 wire _01838_;
 wire _01839_;
 wire _01840_;
 wire _01841_;
 wire _01842_;
 wire _01843_;
 wire _01844_;
 wire _01845_;
 wire _01846_;
 wire _01847_;
 wire _01848_;
 wire _01849_;
 wire _01850_;
 wire _01851_;
 wire _01852_;
 wire _01853_;
 wire _01854_;
 wire _01855_;
 wire _01856_;
 wire _01857_;
 wire _01858_;
 wire _01859_;
 wire _01860_;
 wire _01861_;
 wire _01862_;
 wire _01863_;
 wire _01864_;
 wire _01865_;
 wire _01866_;
 wire _01867_;
 wire _01868_;
 wire _01869_;
 wire _01870_;
 wire _01871_;
 wire _01872_;
 wire _01873_;
 wire _01874_;
 wire _01875_;
 wire _01876_;
 wire _01877_;
 wire _01878_;
 wire _01879_;
 wire _01880_;
 wire _01881_;
 wire _01882_;
 wire _01883_;
 wire _01884_;
 wire _01885_;
 wire _01886_;
 wire _01887_;
 wire _01888_;
 wire _01889_;
 wire _01890_;
 wire _01891_;
 wire _01892_;
 wire _01893_;
 wire _01894_;
 wire _01895_;
 wire _01896_;
 wire _01897_;
 wire _01898_;
 wire _01899_;
 wire _01900_;
 wire _01901_;
 wire _01902_;
 wire _01903_;
 wire _01904_;
 wire _01905_;
 wire _01906_;
 wire _01907_;
 wire _01908_;
 wire _01909_;
 wire _01910_;
 wire _01911_;
 wire _01912_;
 wire _01913_;
 wire _01914_;
 wire _01915_;
 wire _01916_;
 wire _01917_;
 wire _01918_;
 wire _01919_;
 wire _01920_;
 wire _01921_;
 wire _01922_;
 wire _01923_;
 wire _01924_;
 wire _01925_;
 wire _01926_;
 wire _01927_;
 wire _01928_;
 wire _01929_;
 wire _01930_;
 wire _01931_;
 wire _01932_;
 wire _01933_;
 wire _01934_;
 wire _01935_;
 wire _01936_;
 wire _01937_;
 wire _01938_;
 wire _01939_;
 wire _01940_;
 wire _01941_;
 wire _01942_;
 wire _01943_;
 wire _01944_;
 wire _01945_;
 wire _01946_;
 wire _01947_;
 wire _01948_;
 wire _01949_;
 wire _01950_;
 wire _01951_;
 wire _01952_;
 wire _01953_;
 wire _01954_;
 wire _01955_;
 wire _01956_;
 wire _01957_;
 wire _01958_;
 wire _01959_;
 wire _01960_;
 wire _01961_;
 wire _01962_;
 wire _01963_;
 wire _01964_;
 wire _01965_;
 wire _01966_;
 wire _01967_;
 wire _01968_;
 wire _01969_;
 wire _01970_;
 wire _01971_;
 wire _01972_;
 wire _01973_;
 wire _01974_;
 wire _01975_;
 wire _01976_;
 wire _01977_;
 wire _01978_;
 wire _01979_;
 wire _01980_;
 wire _01981_;
 wire _01982_;
 wire _01983_;
 wire _01984_;
 wire _01985_;
 wire _01986_;
 wire _01987_;
 wire _01988_;
 wire _01989_;
 wire _01990_;
 wire _01991_;
 wire _01992_;
 wire _01993_;
 wire _01994_;
 wire _01995_;
 wire _01996_;
 wire _01997_;
 wire _01998_;
 wire _01999_;
 wire _02000_;
 wire _02001_;
 wire _02002_;
 wire _02003_;
 wire _02004_;
 wire _02005_;
 wire _02006_;
 wire _02007_;
 wire _02008_;
 wire _02009_;
 wire _02010_;
 wire _02011_;
 wire _02012_;
 wire _02013_;
 wire _02014_;
 wire _02015_;
 wire _02016_;
 wire _02017_;
 wire _02018_;
 wire _02019_;
 wire _02020_;
 wire _02021_;
 wire _02022_;
 wire _02023_;
 wire _02024_;
 wire _02025_;
 wire _02026_;
 wire _02027_;
 wire _02028_;
 wire _02029_;
 wire _02030_;
 wire _02031_;
 wire _02032_;
 wire _02033_;
 wire _02034_;
 wire _02035_;
 wire _02036_;
 wire _02037_;
 wire _02038_;
 wire _02039_;
 wire _02040_;
 wire _02041_;
 wire _02042_;
 wire _02043_;
 wire _02044_;
 wire _02045_;
 wire _02046_;
 wire _02047_;
 wire _02048_;
 wire _02049_;
 wire _02050_;
 wire _02051_;
 wire _02052_;
 wire _02053_;
 wire _02054_;
 wire _02055_;
 wire _02056_;
 wire _02057_;
 wire _02058_;
 wire _02059_;
 wire _02060_;
 wire _02061_;
 wire _02062_;
 wire _02063_;
 wire _02064_;
 wire _02065_;
 wire _02066_;
 wire _02067_;
 wire _02068_;
 wire _02069_;
 wire _02070_;
 wire _02071_;
 wire _02072_;
 wire _02073_;
 wire _02074_;
 wire _02075_;
 wire _02076_;
 wire _02077_;
 wire _02078_;
 wire _02079_;
 wire _02080_;
 wire _02081_;
 wire _02082_;
 wire _02083_;
 wire _02084_;
 wire _02085_;
 wire _02086_;
 wire _02087_;
 wire _02088_;
 wire _02089_;
 wire _02090_;
 wire _02091_;
 wire _02092_;
 wire _02093_;
 wire _02094_;
 wire _02095_;
 wire _02096_;
 wire _02097_;
 wire _02098_;
 wire _02099_;
 wire _02100_;
 wire _02101_;
 wire _02102_;
 wire _02103_;
 wire _02104_;
 wire _02105_;
 wire _02106_;
 wire _02107_;
 wire _02108_;
 wire _02109_;
 wire _02110_;
 wire _02111_;
 wire _02112_;
 wire _02113_;
 wire _02114_;
 wire _02115_;
 wire _02116_;
 wire _02117_;
 wire _02118_;
 wire _02119_;
 wire _02120_;
 wire _02121_;
 wire _02122_;
 wire _02123_;
 wire _02124_;
 wire _02125_;
 wire _02126_;
 wire _02127_;
 wire _02128_;
 wire _02129_;
 wire _02130_;
 wire _02131_;
 wire _02132_;
 wire _02133_;
 wire _02134_;
 wire _02135_;
 wire _02136_;
 wire _02137_;
 wire _02138_;
 wire _02139_;
 wire _02140_;
 wire _02141_;
 wire _02142_;
 wire _02143_;
 wire _02144_;
 wire _02145_;
 wire _02146_;
 wire _02147_;
 wire _02148_;
 wire _02149_;
 wire _02150_;
 wire _02151_;
 wire _02152_;
 wire _02153_;
 wire _02154_;
 wire _02155_;
 wire _02156_;
 wire _02157_;
 wire _02158_;
 wire _02159_;
 wire _02160_;
 wire _02161_;
 wire _02162_;
 wire _02163_;
 wire _02164_;
 wire _02165_;
 wire _02166_;
 wire _02167_;
 wire _02168_;
 wire _02169_;
 wire _02170_;
 wire _02171_;
 wire _02172_;
 wire _02173_;
 wire _02174_;
 wire _02175_;
 wire _02176_;
 wire _02177_;
 wire _02178_;
 wire _02179_;
 wire _02180_;
 wire _02181_;
 wire _02182_;
 wire _02183_;
 wire _02184_;
 wire _02185_;
 wire _02186_;
 wire _02187_;
 wire _02188_;
 wire _02189_;
 wire _02190_;
 wire _02191_;
 wire _02192_;
 wire _02193_;
 wire _02194_;
 wire _02195_;
 wire _02196_;
 wire _02197_;
 wire _02198_;
 wire _02199_;
 wire _02200_;
 wire _02201_;
 wire _02202_;
 wire _02203_;
 wire _02204_;
 wire _02205_;
 wire _02206_;
 wire _02207_;
 wire _02208_;
 wire _02209_;
 wire _02210_;
 wire _02211_;
 wire _02212_;
 wire _02213_;
 wire _02214_;
 wire _02215_;
 wire _02216_;
 wire _02217_;
 wire _02218_;
 wire _02219_;
 wire _02220_;
 wire _02221_;
 wire _02222_;
 wire _02223_;
 wire _02224_;
 wire _02225_;
 wire _02226_;
 wire _02227_;
 wire _02228_;
 wire _02229_;
 wire _02230_;
 wire _02231_;
 wire _02232_;
 wire _02233_;
 wire _02234_;
 wire _02235_;
 wire _02236_;
 wire _02237_;
 wire _02238_;
 wire _02239_;
 wire _02240_;
 wire _02241_;
 wire _02242_;
 wire _02243_;
 wire _02244_;
 wire _02245_;
 wire _02246_;
 wire _02247_;
 wire _02248_;
 wire _02249_;
 wire _02250_;
 wire _02251_;
 wire _02252_;
 wire _02253_;
 wire _02254_;
 wire _02255_;
 wire _02256_;
 wire _02257_;
 wire _02258_;
 wire _02259_;
 wire _02260_;
 wire _02261_;
 wire _02262_;
 wire _02263_;
 wire _02264_;
 wire _02265_;
 wire _02266_;
 wire _02267_;
 wire _02268_;
 wire _02269_;
 wire _02270_;
 wire _02271_;
 wire _02272_;
 wire _02273_;
 wire _02274_;
 wire _02275_;
 wire _02276_;
 wire _02277_;
 wire _02278_;
 wire _02279_;
 wire _02280_;
 wire _02281_;
 wire _02282_;
 wire _02283_;
 wire _02284_;
 wire _02285_;
 wire _02286_;
 wire _02287_;
 wire _02288_;
 wire _02289_;
 wire _02290_;
 wire _02291_;
 wire _02292_;
 wire _02293_;
 wire _02294_;
 wire _02295_;
 wire _02296_;
 wire _02297_;
 wire _02298_;
 wire _02299_;
 wire _02300_;
 wire _02301_;
 wire _02302_;
 wire _02303_;
 wire _02304_;
 wire _02305_;
 wire _02306_;
 wire _02307_;
 wire _02308_;
 wire _02309_;
 wire _02310_;
 wire _02311_;
 wire _02312_;
 wire _02313_;
 wire _02314_;
 wire _02315_;
 wire _02316_;
 wire _02317_;
 wire _02318_;
 wire _02319_;
 wire _02320_;
 wire _02321_;
 wire _02322_;
 wire _02323_;
 wire _02324_;
 wire _02325_;
 wire _02326_;
 wire _02327_;
 wire _02328_;
 wire _02329_;
 wire _02330_;
 wire _02331_;
 wire _02332_;
 wire _02333_;
 wire _02334_;
 wire _02335_;
 wire _02336_;
 wire _02337_;
 wire _02338_;
 wire _02339_;
 wire _02340_;
 wire _02341_;
 wire _02342_;
 wire _02343_;
 wire _02344_;
 wire _02345_;
 wire _02346_;
 wire _02347_;
 wire _02348_;
 wire _02349_;
 wire _02350_;
 wire _02351_;
 wire _02352_;
 wire _02353_;
 wire _02354_;
 wire _02355_;
 wire _02356_;
 wire _02357_;
 wire _02358_;
 wire _02359_;
 wire _02360_;
 wire _02361_;
 wire _02362_;
 wire _02363_;
 wire _02364_;
 wire _02365_;
 wire _02366_;
 wire _02367_;
 wire _02368_;
 wire _02369_;
 wire _02370_;
 wire _02371_;
 wire _02372_;
 wire _02373_;
 wire _02374_;
 wire _02375_;
 wire _02376_;
 wire _02377_;
 wire _02378_;
 wire _02379_;
 wire _02380_;
 wire _02381_;
 wire _02382_;
 wire _02383_;
 wire _02384_;
 wire _02385_;
 wire _02386_;
 wire _02387_;
 wire _02388_;
 wire _02389_;
 wire _02390_;
 wire _02391_;
 wire _02392_;
 wire _02393_;
 wire _02394_;
 wire _02395_;
 wire _02396_;
 wire _02397_;
 wire _02398_;
 wire _02399_;
 wire _02400_;
 wire _02401_;
 wire _02402_;
 wire _02403_;
 wire _02404_;
 wire _02405_;
 wire _02406_;
 wire _02407_;
 wire _02408_;
 wire _02409_;
 wire _02410_;
 wire _02411_;
 wire _02412_;
 wire _02413_;
 wire _02414_;
 wire _02415_;
 wire _02416_;
 wire _02417_;
 wire _02418_;
 wire _02419_;
 wire _02420_;
 wire _02421_;
 wire _02422_;
 wire _02423_;
 wire _02424_;
 wire _02425_;
 wire _02426_;
 wire _02427_;
 wire _02428_;
 wire _02429_;
 wire _02430_;
 wire _02431_;
 wire _02432_;
 wire _02433_;
 wire _02434_;
 wire _02435_;
 wire _02436_;
 wire _02437_;
 wire _02438_;
 wire _02439_;
 wire _02440_;
 wire _02441_;
 wire _02442_;
 wire _02443_;
 wire _02444_;
 wire _02445_;
 wire _02446_;
 wire _02447_;
 wire _02448_;
 wire _02449_;
 wire _02450_;
 wire _02451_;
 wire _02452_;
 wire _02453_;
 wire _02454_;
 wire _02455_;
 wire _02456_;
 wire _02457_;
 wire _02458_;
 wire _02459_;
 wire _02460_;
 wire _02461_;
 wire _02462_;
 wire _02463_;
 wire _02464_;
 wire _02465_;
 wire _02466_;
 wire _02467_;
 wire _02468_;
 wire _02469_;
 wire _02470_;
 wire _02471_;
 wire _02472_;
 wire _02473_;
 wire _02474_;
 wire _02475_;
 wire _02476_;
 wire _02477_;
 wire _02478_;
 wire _02479_;
 wire _02480_;
 wire _02481_;
 wire _02482_;
 wire _02483_;
 wire _02484_;
 wire _02485_;
 wire _02486_;
 wire _02487_;
 wire _02488_;
 wire _02489_;
 wire _02490_;
 wire _02491_;
 wire _02492_;
 wire _02493_;
 wire _02494_;
 wire _02495_;
 wire _02496_;
 wire _02497_;
 wire _02498_;
 wire _02499_;
 wire _02500_;
 wire _02501_;
 wire _02502_;
 wire _02503_;
 wire _02504_;
 wire _02505_;
 wire _02506_;
 wire _02507_;
 wire _02508_;
 wire _02509_;
 wire _02510_;
 wire _02511_;
 wire _02512_;
 wire _02513_;
 wire _02514_;
 wire _02515_;
 wire _02516_;
 wire _02517_;
 wire _02518_;
 wire _02519_;
 wire _02520_;
 wire _02521_;
 wire _02522_;
 wire _02523_;
 wire _02524_;
 wire _02525_;
 wire _02526_;
 wire _02527_;
 wire _02528_;
 wire _02529_;
 wire _02530_;
 wire _02531_;
 wire _02532_;
 wire _02533_;
 wire _02534_;
 wire _02535_;
 wire _02536_;
 wire _02537_;
 wire _02538_;
 wire _02539_;
 wire _02540_;
 wire _02541_;
 wire _02542_;
 wire _02543_;
 wire _02544_;
 wire _02545_;
 wire _02546_;
 wire _02547_;
 wire _02548_;
 wire _02549_;
 wire _02550_;
 wire _02551_;
 wire _02552_;
 wire _02553_;
 wire _02554_;
 wire _02555_;
 wire _02556_;
 wire _02557_;
 wire _02558_;
 wire _02559_;
 wire _02560_;
 wire _02561_;
 wire _02562_;
 wire _02563_;
 wire _02564_;
 wire _02565_;
 wire _02566_;
 wire _02567_;
 wire _02568_;
 wire _02569_;
 wire _02570_;
 wire _02571_;
 wire _02572_;
 wire _02573_;
 wire _02574_;
 wire _02575_;
 wire _02576_;
 wire _02577_;
 wire _02578_;
 wire _02579_;
 wire _02580_;
 wire _02581_;
 wire _02582_;
 wire _02583_;
 wire _02584_;
 wire _02585_;
 wire _02586_;
 wire _02587_;
 wire _02588_;
 wire _02589_;
 wire _02590_;
 wire _02591_;
 wire _02592_;
 wire _02593_;
 wire _02594_;
 wire _02595_;
 wire _02596_;
 wire _02597_;
 wire _02598_;
 wire _02599_;
 wire _02600_;
 wire _02601_;
 wire _02602_;
 wire _02603_;
 wire _02604_;
 wire _02605_;
 wire _02606_;
 wire _02607_;
 wire _02608_;
 wire _02609_;
 wire _02610_;
 wire _02611_;
 wire _02612_;
 wire _02613_;
 wire _02614_;
 wire _02615_;
 wire _02616_;
 wire _02617_;
 wire _02618_;
 wire _02619_;
 wire _02620_;
 wire _02621_;
 wire _02622_;
 wire _02623_;
 wire _02624_;
 wire _02625_;
 wire _02626_;
 wire _02627_;
 wire _02628_;
 wire _02629_;
 wire _02630_;
 wire _02631_;
 wire _02632_;
 wire _02633_;
 wire _02634_;
 wire _02635_;
 wire _02636_;
 wire _02637_;
 wire _02638_;
 wire _02639_;
 wire _02640_;
 wire _02641_;
 wire _02642_;
 wire _02643_;
 wire _02644_;
 wire _02645_;
 wire _02646_;
 wire _02647_;
 wire _02648_;
 wire _02649_;
 wire _02650_;
 wire _02651_;
 wire _02652_;
 wire _02653_;
 wire _02654_;
 wire _02655_;
 wire _02656_;
 wire _02657_;
 wire _02658_;
 wire _02659_;
 wire _02660_;
 wire _02661_;
 wire _02662_;
 wire _02663_;
 wire _02664_;
 wire _02665_;
 wire _02666_;
 wire _02667_;
 wire _02668_;
 wire _02669_;
 wire _02670_;
 wire _02671_;
 wire _02672_;
 wire _02673_;
 wire _02674_;
 wire _02675_;
 wire _02676_;
 wire _02677_;
 wire _02678_;
 wire _02679_;
 wire _02680_;
 wire _02681_;
 wire _02682_;
 wire _02683_;
 wire _02684_;
 wire _02685_;
 wire _02686_;
 wire _02687_;
 wire _02688_;
 wire _02689_;
 wire _02690_;
 wire _02691_;
 wire _02692_;
 wire _02693_;
 wire _02694_;
 wire _02695_;
 wire _02696_;
 wire _02697_;
 wire _02698_;
 wire _02699_;
 wire _02700_;
 wire _02701_;
 wire _02702_;
 wire _02703_;
 wire _02704_;
 wire _02705_;
 wire _02706_;
 wire _02707_;
 wire _02708_;
 wire _02709_;
 wire _02710_;
 wire _02711_;
 wire _02712_;
 wire _02713_;
 wire _02714_;
 wire _02715_;
 wire _02716_;
 wire _02717_;
 wire _02718_;
 wire _02719_;
 wire _02720_;
 wire _02721_;
 wire _02722_;
 wire _02723_;
 wire _02724_;
 wire _02725_;
 wire _02726_;
 wire _02727_;
 wire _02728_;
 wire _02729_;
 wire _02730_;
 wire _02731_;
 wire _02732_;
 wire _02733_;
 wire _02734_;
 wire _02735_;
 wire _02736_;
 wire _02737_;
 wire _02738_;
 wire _02739_;
 wire _02740_;
 wire _02741_;
 wire _02742_;
 wire _02743_;
 wire _02744_;
 wire _02745_;
 wire _02746_;
 wire _02747_;
 wire _02748_;
 wire _02749_;
 wire _02750_;
 wire _02751_;
 wire _02752_;
 wire _02753_;
 wire _02754_;
 wire _02755_;
 wire _02756_;
 wire _02757_;
 wire _02758_;
 wire _02759_;
 wire _02760_;
 wire _02761_;
 wire _02762_;
 wire _02763_;
 wire _02764_;
 wire _02765_;
 wire _02766_;
 wire _02767_;
 wire _02768_;
 wire _02769_;
 wire _02770_;
 wire _02771_;
 wire _02772_;
 wire _02773_;
 wire _02774_;
 wire _02775_;
 wire _02776_;
 wire _02777_;
 wire _02778_;
 wire _02779_;
 wire _02780_;
 wire _02781_;
 wire _02782_;
 wire _02783_;
 wire _02784_;
 wire _02785_;
 wire _02786_;
 wire _02787_;
 wire _02788_;
 wire _02789_;
 wire _02790_;
 wire _02791_;
 wire _02792_;
 wire _02793_;
 wire _02794_;
 wire _02795_;
 wire _02796_;
 wire _02797_;
 wire _02798_;
 wire _02799_;
 wire _02800_;
 wire _02801_;
 wire _02802_;
 wire _02803_;
 wire _02804_;
 wire _02805_;
 wire _02806_;
 wire _02807_;
 wire _02808_;
 wire _02809_;
 wire _02810_;
 wire _02811_;
 wire _02812_;
 wire _02813_;
 wire _02814_;
 wire _02815_;
 wire _02816_;
 wire _02817_;
 wire _02818_;
 wire _02819_;
 wire _02820_;
 wire _02821_;
 wire _02822_;
 wire _02823_;
 wire _02824_;
 wire _02825_;
 wire _02826_;
 wire _02827_;
 wire _02828_;
 wire _02829_;
 wire _02830_;
 wire _02831_;
 wire _02832_;
 wire _02833_;
 wire _02834_;
 wire _02835_;
 wire _02836_;
 wire _02837_;
 wire _02838_;
 wire _02839_;
 wire _02840_;
 wire _02841_;
 wire _02842_;
 wire _02843_;
 wire _02844_;
 wire _02845_;
 wire _02846_;
 wire _02847_;
 wire _02848_;
 wire _02849_;
 wire _02850_;
 wire _02851_;
 wire _02852_;
 wire _02853_;
 wire _02854_;
 wire _02855_;
 wire _02856_;
 wire _02857_;
 wire _02858_;
 wire _02859_;
 wire _02860_;
 wire _02861_;
 wire _02862_;
 wire _02863_;
 wire _02864_;
 wire _02865_;
 wire _02866_;
 wire _02867_;
 wire _02868_;
 wire _02869_;
 wire _02870_;
 wire _02871_;
 wire _02872_;
 wire _02873_;
 wire _02874_;
 wire _02875_;
 wire _02876_;
 wire _02877_;
 wire _02878_;
 wire _02879_;
 wire _02880_;
 wire _02881_;
 wire _02882_;
 wire _02883_;
 wire _02884_;
 wire _02885_;
 wire _02886_;
 wire _02887_;
 wire _02888_;
 wire _02889_;
 wire _02890_;
 wire _02891_;
 wire _02892_;
 wire _02893_;
 wire _02894_;
 wire _02895_;
 wire _02896_;
 wire _02897_;
 wire _02898_;
 wire _02899_;
 wire _02900_;
 wire _02901_;
 wire _02902_;
 wire _02903_;
 wire _02904_;
 wire _02905_;
 wire _02906_;
 wire _02907_;
 wire _02908_;
 wire _02909_;
 wire _02910_;
 wire _02911_;
 wire _02912_;
 wire _02913_;
 wire _02914_;
 wire _02915_;
 wire _02916_;
 wire _02917_;
 wire _02918_;
 wire _02919_;
 wire _02920_;
 wire _02921_;
 wire _02922_;
 wire _02923_;
 wire _02924_;
 wire _02925_;
 wire _02926_;
 wire _02927_;
 wire _02928_;
 wire _02929_;
 wire _02930_;
 wire _02931_;
 wire _02932_;
 wire _02933_;
 wire _02934_;
 wire _02935_;
 wire _02936_;
 wire _02937_;
 wire _02938_;
 wire _02939_;
 wire _02940_;
 wire _02941_;
 wire _02942_;
 wire _02943_;
 wire _02944_;
 wire _02945_;
 wire _02946_;
 wire _02947_;
 wire _02948_;
 wire _02949_;
 wire _02950_;
 wire _02951_;
 wire _02952_;
 wire _02953_;
 wire _02954_;
 wire _02955_;
 wire _02956_;
 wire _02957_;
 wire _02958_;
 wire _02959_;
 wire _02960_;
 wire _02961_;
 wire _02962_;
 wire _02963_;
 wire _02964_;
 wire _02965_;
 wire _02966_;
 wire _02967_;
 wire _02968_;
 wire _02969_;
 wire _02970_;
 wire _02971_;
 wire _02972_;
 wire _02973_;
 wire _02974_;
 wire _02975_;
 wire _02976_;
 wire _02977_;
 wire _02978_;
 wire _02979_;
 wire _02980_;
 wire _02981_;
 wire _02982_;
 wire _02983_;
 wire _02984_;
 wire _02985_;
 wire _02986_;
 wire _02987_;
 wire _02988_;
 wire _02989_;
 wire _02990_;
 wire _02991_;
 wire _02992_;
 wire _02993_;
 wire _02994_;
 wire _02995_;
 wire _02996_;
 wire _02997_;
 wire _02998_;
 wire _02999_;
 wire _03000_;
 wire _03001_;
 wire _03002_;
 wire _03003_;
 wire _03004_;
 wire _03005_;
 wire _03006_;
 wire _03007_;
 wire _03008_;
 wire _03009_;
 wire _03010_;
 wire _03011_;
 wire _03012_;
 wire _03013_;
 wire _03014_;
 wire _03015_;
 wire _03016_;
 wire _03017_;
 wire _03018_;
 wire _03019_;
 wire _03020_;
 wire _03021_;
 wire _03022_;
 wire _03023_;
 wire _03024_;
 wire _03025_;
 wire _03026_;
 wire _03027_;
 wire _03028_;
 wire _03029_;
 wire _03030_;
 wire _03031_;
 wire _03032_;
 wire _03033_;
 wire _03034_;
 wire _03035_;
 wire _03036_;
 wire _03037_;
 wire _03038_;
 wire _03039_;
 wire _03040_;
 wire _03041_;
 wire _03042_;
 wire _03043_;
 wire _03044_;
 wire _03045_;
 wire _03046_;
 wire _03047_;
 wire _03048_;
 wire _03049_;
 wire _03050_;
 wire _03051_;
 wire _03052_;
 wire _03053_;
 wire _03054_;
 wire _03055_;
 wire _03056_;
 wire _03057_;
 wire _03058_;
 wire _03059_;
 wire _03060_;
 wire _03061_;
 wire _03062_;
 wire _03063_;
 wire _03064_;
 wire _03065_;
 wire _03066_;
 wire _03067_;
 wire _03068_;
 wire _03069_;
 wire _03070_;
 wire _03071_;
 wire _03072_;
 wire _03073_;
 wire _03074_;
 wire _03075_;
 wire _03076_;
 wire _03077_;
 wire _03078_;
 wire _03079_;
 wire _03080_;
 wire _03081_;
 wire _03082_;
 wire _03083_;
 wire _03084_;
 wire _03085_;
 wire _03086_;
 wire _03087_;
 wire _03088_;
 wire _03089_;
 wire _03090_;
 wire _03091_;
 wire _03092_;
 wire _03093_;
 wire _03094_;
 wire _03095_;
 wire _03096_;
 wire _03097_;
 wire _03098_;
 wire _03099_;
 wire _03100_;
 wire _03101_;
 wire _03102_;
 wire _03103_;
 wire _03104_;
 wire _03105_;
 wire _03106_;
 wire _03107_;
 wire _03108_;
 wire _03109_;
 wire _03110_;
 wire _03111_;
 wire _03112_;
 wire _03113_;
 wire _03114_;
 wire _03115_;
 wire _03116_;
 wire _03117_;
 wire _03118_;
 wire _03119_;
 wire _03120_;
 wire _03121_;
 wire _03122_;
 wire _03123_;
 wire _03124_;
 wire _03125_;
 wire _03126_;
 wire _03127_;
 wire _03128_;
 wire _03129_;
 wire _03130_;
 wire _03131_;
 wire _03132_;
 wire _03133_;
 wire _03134_;
 wire _03135_;
 wire _03136_;
 wire _03137_;
 wire _03138_;
 wire _03139_;
 wire _03140_;
 wire _03141_;
 wire _03142_;
 wire _03143_;
 wire _03144_;
 wire _03145_;
 wire _03146_;
 wire _03147_;
 wire _03148_;
 wire _03149_;
 wire _03150_;
 wire _03151_;
 wire _03152_;
 wire _03153_;
 wire _03154_;
 wire _03155_;
 wire _03156_;
 wire _03157_;
 wire _03158_;
 wire _03159_;
 wire _03160_;
 wire _03161_;
 wire _03162_;
 wire _03163_;
 wire _03164_;
 wire _03165_;
 wire _03166_;
 wire _03167_;
 wire _03168_;
 wire _03169_;
 wire _03170_;
 wire _03171_;
 wire _03172_;
 wire _03173_;
 wire _03174_;
 wire _03175_;
 wire _03176_;
 wire _03177_;
 wire _03178_;
 wire _03179_;
 wire _03180_;
 wire _03181_;
 wire _03182_;
 wire _03183_;
 wire _03184_;
 wire _03185_;
 wire _03186_;
 wire _03187_;
 wire _03188_;
 wire _03189_;
 wire _03190_;
 wire _03191_;
 wire _03192_;
 wire _03193_;
 wire _03194_;
 wire _03195_;
 wire _03196_;
 wire _03197_;
 wire _03198_;
 wire _03199_;
 wire _03200_;
 wire _03201_;
 wire _03202_;
 wire _03203_;
 wire _03204_;
 wire _03205_;
 wire _03206_;
 wire _03207_;
 wire _03208_;
 wire _03209_;
 wire _03210_;
 wire _03211_;
 wire _03212_;
 wire _03213_;
 wire _03214_;
 wire _03215_;
 wire _03216_;
 wire _03217_;
 wire _03218_;
 wire _03219_;
 wire _03220_;
 wire _03221_;
 wire _03222_;
 wire _03223_;
 wire _03224_;
 wire _03225_;
 wire _03226_;
 wire _03227_;
 wire _03228_;
 wire _03229_;
 wire _03230_;
 wire _03231_;
 wire _03232_;
 wire _03233_;
 wire _03234_;
 wire _03235_;
 wire _03236_;
 wire _03237_;
 wire _03238_;
 wire _03239_;
 wire _03240_;
 wire _03241_;
 wire _03242_;
 wire _03243_;
 wire _03244_;
 wire _03245_;
 wire _03246_;
 wire _03247_;
 wire _03248_;
 wire _03249_;
 wire _03250_;
 wire _03251_;
 wire _03252_;
 wire _03253_;
 wire _03254_;
 wire _03255_;
 wire _03256_;
 wire _03257_;
 wire _03258_;
 wire _03259_;
 wire _03260_;
 wire _03261_;
 wire _03262_;
 wire _03263_;
 wire _03264_;
 wire _03265_;
 wire _03266_;
 wire _03267_;
 wire _03268_;
 wire _03269_;
 wire _03270_;
 wire _03271_;
 wire _03272_;
 wire _03273_;
 wire _03274_;
 wire _03275_;
 wire _03276_;
 wire _03277_;
 wire _03278_;
 wire _03279_;
 wire _03280_;
 wire _03281_;
 wire _03282_;
 wire _03283_;
 wire _03284_;
 wire _03285_;
 wire _03286_;
 wire _03287_;
 wire _03288_;
 wire _03289_;
 wire _03290_;
 wire _03291_;
 wire _03292_;
 wire _03293_;
 wire _03294_;
 wire _03295_;
 wire _03296_;
 wire _03297_;
 wire _03298_;
 wire _03299_;
 wire _03300_;
 wire _03301_;
 wire _03302_;
 wire _03303_;
 wire _03304_;
 wire _03305_;
 wire _03306_;
 wire _03307_;
 wire _03308_;
 wire _03309_;
 wire _03310_;
 wire _03311_;
 wire _03312_;
 wire _03313_;
 wire _03314_;
 wire _03315_;
 wire _03316_;
 wire _03317_;
 wire _03318_;
 wire _03319_;
 wire _03320_;
 wire _03321_;
 wire _03322_;
 wire _03323_;
 wire _03324_;
 wire _03325_;
 wire _03326_;
 wire _03327_;
 wire _03328_;
 wire _03329_;
 wire _03330_;
 wire _03331_;
 wire _03332_;
 wire _03333_;
 wire _03334_;
 wire _03335_;
 wire _03336_;
 wire _03337_;
 wire _03338_;
 wire _03339_;
 wire _03340_;
 wire _03341_;
 wire _03342_;
 wire _03343_;
 wire _03344_;
 wire _03345_;
 wire _03346_;
 wire _03347_;
 wire _03348_;
 wire _03349_;
 wire _03350_;
 wire _03351_;
 wire _03352_;
 wire _03353_;
 wire _03354_;
 wire _03355_;
 wire _03356_;
 wire _03357_;
 wire _03358_;
 wire _03359_;
 wire _03360_;
 wire _03361_;
 wire _03362_;
 wire _03363_;
 wire _03364_;
 wire _03365_;
 wire _03366_;
 wire _03367_;
 wire _03368_;
 wire _03369_;
 wire _03370_;
 wire _03371_;
 wire _03372_;
 wire _03373_;
 wire _03374_;
 wire _03375_;
 wire _03376_;
 wire _03377_;
 wire _03378_;
 wire _03379_;
 wire _03380_;
 wire _03381_;
 wire _03382_;
 wire _03383_;
 wire _03384_;
 wire _03385_;
 wire _03386_;
 wire _03387_;
 wire _03388_;
 wire _03389_;
 wire _03390_;
 wire _03391_;
 wire _03392_;
 wire _03393_;
 wire _03394_;
 wire _03395_;
 wire _03396_;
 wire _03397_;
 wire _03398_;
 wire _03399_;
 wire _03400_;
 wire _03401_;
 wire _03402_;
 wire _03403_;
 wire _03404_;
 wire _03405_;
 wire _03406_;
 wire _03407_;
 wire _03408_;
 wire _03409_;
 wire _03410_;
 wire _03411_;
 wire _03412_;
 wire _03413_;
 wire _03414_;
 wire _03415_;
 wire _03416_;
 wire _03417_;
 wire _03418_;
 wire _03419_;
 wire _03420_;
 wire _03421_;
 wire _03422_;
 wire _03423_;
 wire _03424_;
 wire _03425_;
 wire _03426_;
 wire _03427_;
 wire _03428_;
 wire _03429_;
 wire _03430_;
 wire _03431_;
 wire _03432_;
 wire _03433_;
 wire _03434_;
 wire _03435_;
 wire _03436_;
 wire _03437_;
 wire _03438_;
 wire _03439_;
 wire _03440_;
 wire _03441_;
 wire _03442_;
 wire _03443_;
 wire _03444_;
 wire _03445_;
 wire _03446_;
 wire _03447_;
 wire _03448_;
 wire _03449_;
 wire _03450_;
 wire _03451_;
 wire _03452_;
 wire _03453_;
 wire _03454_;
 wire _03455_;
 wire _03456_;
 wire _03457_;
 wire _03458_;
 wire _03459_;
 wire _03460_;
 wire _03461_;
 wire _03462_;
 wire _03463_;
 wire _03464_;
 wire _03465_;
 wire _03466_;
 wire _03467_;
 wire _03468_;
 wire _03469_;
 wire _03470_;
 wire _03471_;
 wire _03472_;
 wire _03473_;
 wire _03474_;
 wire _03475_;
 wire _03476_;
 wire _03477_;
 wire _03478_;
 wire _03479_;
 wire _03480_;
 wire _03481_;
 wire _03482_;
 wire _03483_;
 wire _03484_;
 wire _03485_;
 wire _03486_;
 wire _03487_;
 wire _03488_;
 wire _03489_;
 wire _03490_;
 wire _03491_;
 wire _03492_;
 wire _03493_;
 wire _03494_;
 wire _03495_;
 wire _03496_;
 wire _03497_;
 wire _03498_;
 wire _03499_;
 wire _03500_;
 wire _03501_;
 wire _03502_;
 wire _03503_;
 wire _03504_;
 wire _03505_;
 wire _03506_;
 wire _03507_;
 wire _03508_;
 wire _03509_;
 wire _03510_;
 wire _03511_;
 wire _03512_;
 wire _03513_;
 wire _03514_;
 wire _03515_;
 wire _03516_;
 wire _03517_;
 wire _03518_;
 wire _03519_;
 wire _03520_;
 wire _03521_;
 wire _03522_;
 wire _03523_;
 wire _03524_;
 wire _03525_;
 wire _03526_;
 wire _03527_;
 wire _03528_;
 wire _03529_;
 wire _03530_;
 wire _03531_;
 wire _03532_;
 wire _03533_;
 wire _03534_;
 wire _03535_;
 wire _03536_;
 wire _03537_;
 wire _03538_;
 wire _03539_;
 wire _03540_;
 wire _03541_;
 wire _03542_;
 wire _03543_;
 wire _03544_;
 wire _03545_;
 wire _03546_;
 wire _03547_;
 wire _03548_;
 wire _03549_;
 wire _03550_;
 wire _03551_;
 wire _03552_;
 wire _03553_;
 wire _03554_;
 wire _03555_;
 wire _03556_;
 wire _03557_;
 wire _03558_;
 wire _03559_;
 wire _03560_;
 wire _03561_;
 wire _03562_;
 wire _03563_;
 wire _03564_;
 wire _03565_;
 wire _03566_;
 wire _03567_;
 wire _03568_;
 wire _03569_;
 wire _03570_;
 wire _03571_;
 wire _03572_;
 wire _03573_;
 wire _03574_;
 wire _03575_;
 wire _03576_;
 wire _03577_;
 wire _03578_;
 wire _03579_;
 wire _03580_;
 wire _03581_;
 wire _03582_;
 wire _03583_;
 wire _03584_;
 wire _03585_;
 wire _03586_;
 wire _03587_;
 wire _03588_;
 wire _03589_;
 wire _03590_;
 wire _03591_;
 wire _03592_;
 wire _03593_;
 wire _03594_;
 wire _03595_;
 wire _03596_;
 wire _03597_;
 wire _03598_;
 wire _03599_;
 wire _03600_;
 wire _03601_;
 wire _03602_;
 wire _03603_;
 wire _03604_;
 wire _03605_;
 wire _03606_;
 wire _03607_;
 wire _03608_;
 wire _03609_;
 wire _03610_;
 wire _03611_;
 wire _03612_;
 wire _03613_;
 wire _03614_;
 wire _03615_;
 wire _03616_;
 wire _03617_;
 wire _03618_;
 wire _03619_;
 wire _03620_;
 wire _03621_;
 wire _03622_;
 wire _03623_;
 wire _03624_;
 wire _03625_;
 wire _03626_;
 wire _03627_;
 wire _03628_;
 wire _03629_;
 wire _03630_;
 wire _03631_;
 wire _03632_;
 wire _03633_;
 wire _03634_;
 wire _03635_;
 wire _03636_;
 wire _03637_;
 wire _03638_;
 wire _03639_;
 wire _03640_;
 wire _03641_;
 wire _03642_;
 wire _03643_;
 wire _03644_;
 wire _03645_;
 wire _03646_;
 wire _03647_;
 wire _03648_;
 wire _03649_;
 wire _03650_;
 wire _03651_;
 wire _03652_;
 wire _03653_;
 wire _03654_;
 wire _03655_;
 wire _03656_;
 wire _03657_;
 wire _03658_;
 wire _03659_;
 wire _03660_;
 wire _03661_;
 wire _03662_;
 wire _03663_;
 wire _03664_;
 wire _03665_;
 wire _03666_;
 wire _03667_;
 wire _03668_;
 wire _03669_;
 wire _03670_;
 wire _03671_;
 wire _03672_;
 wire _03673_;
 wire _03674_;
 wire _03675_;
 wire _03676_;
 wire _03677_;
 wire _03678_;
 wire _03679_;
 wire _03680_;
 wire _03681_;
 wire _03682_;
 wire _03683_;
 wire _03684_;
 wire _03685_;
 wire _03686_;
 wire _03687_;
 wire _03688_;
 wire _03689_;
 wire _03690_;
 wire _03691_;
 wire _03692_;
 wire _03693_;
 wire _03694_;
 wire _03695_;
 wire _03696_;
 wire _03697_;
 wire _03698_;
 wire _03699_;
 wire _03700_;
 wire _03701_;
 wire _03702_;
 wire _03703_;
 wire _03704_;
 wire _03705_;
 wire _03706_;
 wire _03707_;
 wire _03708_;
 wire _03709_;
 wire _03710_;
 wire _03711_;
 wire _03712_;
 wire _03713_;
 wire _03714_;
 wire _03715_;
 wire _03716_;
 wire _03717_;
 wire _03718_;
 wire _03719_;
 wire _03720_;
 wire _03721_;
 wire _03722_;
 wire _03723_;
 wire _03724_;
 wire _03725_;
 wire _03726_;
 wire _03727_;
 wire _03728_;
 wire _03729_;
 wire _03730_;
 wire _03731_;
 wire _03732_;
 wire _03733_;
 wire _03734_;
 wire _03735_;
 wire _03736_;
 wire _03737_;
 wire _03738_;
 wire _03739_;
 wire _03740_;
 wire _03741_;
 wire _03742_;
 wire _03743_;
 wire _03744_;
 wire _03745_;
 wire _03746_;
 wire _03747_;
 wire _03748_;
 wire _03749_;
 wire _03750_;
 wire _03751_;
 wire _03752_;
 wire _03753_;
 wire _03754_;
 wire _03755_;
 wire _03756_;
 wire _03757_;
 wire _03758_;
 wire _03759_;
 wire _03760_;
 wire _03761_;
 wire _03762_;
 wire _03763_;
 wire _03764_;
 wire _03765_;
 wire _03766_;
 wire _03767_;
 wire _03768_;
 wire _03769_;
 wire _03770_;
 wire _03771_;
 wire _03772_;
 wire _03773_;
 wire _03774_;
 wire _03775_;
 wire _03776_;
 wire _03777_;
 wire _03778_;
 wire _03779_;
 wire _03780_;
 wire _03781_;
 wire _03782_;
 wire _03783_;
 wire _03784_;
 wire _03785_;
 wire _03786_;
 wire _03787_;
 wire _03788_;
 wire _03789_;
 wire _03790_;
 wire _03791_;
 wire _03792_;
 wire _03793_;
 wire _03794_;
 wire _03795_;
 wire _03796_;
 wire _03797_;
 wire _03798_;
 wire _03799_;
 wire _03800_;
 wire _03801_;
 wire _03802_;
 wire _03803_;
 wire _03804_;
 wire _03805_;
 wire _03806_;
 wire _03807_;
 wire _03808_;
 wire _03809_;
 wire _03810_;
 wire _03811_;
 wire _03812_;
 wire _03813_;
 wire _03814_;
 wire _03815_;
 wire _03816_;
 wire _03817_;
 wire _03818_;
 wire _03819_;
 wire _03820_;
 wire _03821_;
 wire _03822_;
 wire _03823_;
 wire _03824_;
 wire _03825_;
 wire _03826_;
 wire _03827_;
 wire _03828_;
 wire _03829_;
 wire _03830_;
 wire _03831_;
 wire _03832_;
 wire _03833_;
 wire _03834_;
 wire _03835_;
 wire _03836_;
 wire _03837_;
 wire _03838_;
 wire _03839_;
 wire _03840_;
 wire _03841_;
 wire _03842_;
 wire _03843_;
 wire _03844_;
 wire _03845_;
 wire _03846_;
 wire _03847_;
 wire _03848_;
 wire _03849_;
 wire _03850_;
 wire _03851_;
 wire _03852_;
 wire _03853_;
 wire _03854_;
 wire _03855_;
 wire _03856_;
 wire _03857_;
 wire _03858_;
 wire _03859_;
 wire _03860_;
 wire _03861_;
 wire _03862_;
 wire _03863_;
 wire _03864_;
 wire _03865_;
 wire _03866_;
 wire _03867_;
 wire _03868_;
 wire _03869_;
 wire _03870_;
 wire _03871_;
 wire _03872_;
 wire _03873_;
 wire _03874_;
 wire _03875_;
 wire _03876_;
 wire _03877_;
 wire _03878_;
 wire _03879_;
 wire _03880_;
 wire _03881_;
 wire _03882_;
 wire _03883_;
 wire _03884_;
 wire _03885_;
 wire _03886_;
 wire _03887_;
 wire _03888_;
 wire _03889_;
 wire _03890_;
 wire _03891_;
 wire _03892_;
 wire _03893_;
 wire _03894_;
 wire _03895_;
 wire _03896_;
 wire _03897_;
 wire _03898_;
 wire _03899_;
 wire _03900_;
 wire _03901_;
 wire _03902_;
 wire _03903_;
 wire _03904_;
 wire _03905_;
 wire _03906_;
 wire _03907_;
 wire _03908_;
 wire _03909_;
 wire _03910_;
 wire _03911_;
 wire _03912_;
 wire _03913_;
 wire _03914_;
 wire _03915_;
 wire _03916_;
 wire _03917_;
 wire _03918_;
 wire _03919_;
 wire _03920_;
 wire _03921_;
 wire _03922_;
 wire _03923_;
 wire _03924_;
 wire _03925_;
 wire _03926_;
 wire _03927_;
 wire _03928_;
 wire _03929_;
 wire _03930_;
 wire _03931_;
 wire _03932_;
 wire _03933_;
 wire _03934_;
 wire _03935_;
 wire _03936_;
 wire _03937_;
 wire _03938_;
 wire _03939_;
 wire _03940_;
 wire _03941_;
 wire _03942_;
 wire _03943_;
 wire _03944_;
 wire _03945_;
 wire _03946_;
 wire _03947_;
 wire _03948_;
 wire _03949_;
 wire _03950_;
 wire _03951_;
 wire _03952_;
 wire _03953_;
 wire _03954_;
 wire _03955_;
 wire _03956_;
 wire _03957_;
 wire _03958_;
 wire _03959_;
 wire _03960_;
 wire _03961_;
 wire _03962_;
 wire _03963_;
 wire _03964_;
 wire _03965_;
 wire _03966_;
 wire _03967_;
 wire _03968_;
 wire _03969_;
 wire _03970_;
 wire _03971_;
 wire _03972_;
 wire _03973_;
 wire _03974_;
 wire _03975_;
 wire _03976_;
 wire _03977_;
 wire _03978_;
 wire _03979_;
 wire _03980_;
 wire _03981_;
 wire _03982_;
 wire _03983_;
 wire _03984_;
 wire _03985_;
 wire _03986_;
 wire _03987_;
 wire _03988_;
 wire _03989_;
 wire _03990_;
 wire _03991_;
 wire _03992_;
 wire _03993_;
 wire _03994_;
 wire _03995_;
 wire _03996_;
 wire _03997_;
 wire _03998_;
 wire _03999_;
 wire _04000_;
 wire _04001_;
 wire _04002_;
 wire _04003_;
 wire _04004_;
 wire _04005_;
 wire _04006_;
 wire _04007_;
 wire _04008_;
 wire _04009_;
 wire _04010_;
 wire _04011_;
 wire _04012_;
 wire _04013_;
 wire _04014_;
 wire _04015_;
 wire _04016_;
 wire _04017_;
 wire _04018_;
 wire _04019_;
 wire _04020_;
 wire _04021_;
 wire _04022_;
 wire _04023_;
 wire _04024_;
 wire _04025_;
 wire _04026_;
 wire _04027_;
 wire _04028_;
 wire _04029_;
 wire _04030_;
 wire _04031_;
 wire _04032_;
 wire _04033_;
 wire _04034_;
 wire _04035_;
 wire _04036_;
 wire _04037_;
 wire _04038_;
 wire _04039_;
 wire _04040_;
 wire _04041_;
 wire _04042_;
 wire _04043_;
 wire _04044_;
 wire _04045_;
 wire _04046_;
 wire _04047_;
 wire _04048_;
 wire _04049_;
 wire _04050_;
 wire _04051_;
 wire _04052_;
 wire _04053_;
 wire _04054_;
 wire _04055_;
 wire _04056_;
 wire _04057_;
 wire _04058_;
 wire _04059_;
 wire _04060_;
 wire _04061_;
 wire _04062_;
 wire _04063_;
 wire _04064_;
 wire _04065_;
 wire _04066_;
 wire _04067_;
 wire _04068_;
 wire _04069_;
 wire _04070_;
 wire _04071_;
 wire _04072_;
 wire _04073_;
 wire _04074_;
 wire _04075_;
 wire _04076_;
 wire _04077_;
 wire _04078_;
 wire _04079_;
 wire _04080_;
 wire _04081_;
 wire _04082_;
 wire _04083_;
 wire _04084_;
 wire _04085_;
 wire _04086_;
 wire _04087_;
 wire _04088_;
 wire _04089_;
 wire _04090_;
 wire _04091_;
 wire _04092_;
 wire _04093_;
 wire _04094_;
 wire _04095_;
 wire _04096_;
 wire _04097_;
 wire _04098_;
 wire _04099_;
 wire _04100_;
 wire _04101_;
 wire _04102_;
 wire _04103_;
 wire _04104_;
 wire _04105_;
 wire _04106_;
 wire _04107_;
 wire _04108_;
 wire _04109_;
 wire _04110_;
 wire _04111_;
 wire _04112_;
 wire _04113_;
 wire _04114_;
 wire _04115_;
 wire _04116_;
 wire _04117_;
 wire _04118_;
 wire _04119_;
 wire _04120_;
 wire _04121_;
 wire _04122_;
 wire _04123_;
 wire _04124_;
 wire _04125_;
 wire _04126_;
 wire _04127_;
 wire _04128_;
 wire _04129_;
 wire _04130_;
 wire _04131_;
 wire _04132_;
 wire _04133_;
 wire _04134_;
 wire _04135_;
 wire _04136_;
 wire _04137_;
 wire _04138_;
 wire _04139_;
 wire _04140_;
 wire _04141_;
 wire _04142_;
 wire _04143_;
 wire _04144_;
 wire _04145_;
 wire _04146_;
 wire _04147_;
 wire _04148_;
 wire _04149_;
 wire _04150_;
 wire _04151_;
 wire _04152_;
 wire _04153_;
 wire _04154_;
 wire _04155_;
 wire _04156_;
 wire _04157_;
 wire _04158_;
 wire _04159_;
 wire _04160_;
 wire _04161_;
 wire _04162_;
 wire _04163_;
 wire _04164_;
 wire _04165_;
 wire _04166_;
 wire _04167_;
 wire _04168_;
 wire _04169_;
 wire _04170_;
 wire _04171_;
 wire _04172_;
 wire _04173_;
 wire _04174_;
 wire _04175_;
 wire _04176_;
 wire _04177_;
 wire _04178_;
 wire _04179_;
 wire _04180_;
 wire _04181_;
 wire _04182_;
 wire _04183_;
 wire _04184_;
 wire _04185_;
 wire _04186_;
 wire _04187_;
 wire _04188_;
 wire _04189_;
 wire _04190_;
 wire _04191_;
 wire _04192_;
 wire _04193_;
 wire _04194_;
 wire _04195_;
 wire _04196_;
 wire _04197_;
 wire _04198_;
 wire _04199_;
 wire _04200_;
 wire _04201_;
 wire _04202_;
 wire _04203_;
 wire _04204_;
 wire _04205_;
 wire _04206_;
 wire _04207_;
 wire _04208_;
 wire _04209_;
 wire _04210_;
 wire _04211_;
 wire _04212_;
 wire _04213_;
 wire _04214_;
 wire _04215_;
 wire _04216_;
 wire _04217_;
 wire _04218_;
 wire _04219_;
 wire _04220_;
 wire _04221_;
 wire _04222_;
 wire _04223_;
 wire _04224_;
 wire _04225_;
 wire _04226_;
 wire _04227_;
 wire _04228_;
 wire _04229_;
 wire _04230_;
 wire _04231_;
 wire _04232_;
 wire _04233_;
 wire _04234_;
 wire _04235_;
 wire _04236_;
 wire _04237_;
 wire _04238_;
 wire _04239_;
 wire _04240_;
 wire _04241_;
 wire _04242_;
 wire _04243_;
 wire _04244_;
 wire _04245_;
 wire _04246_;
 wire _04247_;
 wire _04248_;
 wire _04249_;
 wire _04250_;
 wire _04251_;
 wire _04252_;
 wire _04253_;
 wire _04254_;
 wire _04255_;
 wire _04256_;
 wire _04257_;
 wire _04258_;
 wire _04259_;
 wire _04260_;
 wire _04261_;
 wire _04262_;
 wire _04263_;
 wire _04264_;
 wire _04265_;
 wire _04266_;
 wire _04267_;
 wire _04268_;
 wire _04269_;
 wire _04270_;
 wire _04271_;
 wire _04272_;
 wire _04273_;
 wire _04274_;
 wire _04275_;
 wire _04276_;
 wire _04277_;
 wire _04278_;
 wire _04279_;
 wire _04280_;
 wire _04281_;
 wire _04282_;
 wire _04283_;
 wire _04284_;
 wire _04285_;
 wire _04286_;
 wire _04287_;
 wire _04288_;
 wire _04289_;
 wire _04290_;
 wire _04291_;
 wire _04292_;
 wire _04293_;
 wire _04294_;
 wire _04295_;
 wire _04296_;
 wire _04297_;
 wire _04298_;
 wire _04299_;
 wire _04300_;
 wire _04301_;
 wire _04302_;
 wire _04303_;
 wire _04304_;
 wire _04305_;
 wire _04306_;
 wire _04307_;
 wire _04308_;
 wire _04309_;
 wire _04310_;
 wire _04311_;
 wire _04312_;
 wire _04313_;
 wire _04314_;
 wire _04315_;
 wire _04316_;
 wire _04317_;
 wire _04318_;
 wire _04319_;
 wire _04320_;
 wire _04321_;
 wire _04322_;
 wire _04323_;
 wire _04324_;
 wire _04325_;
 wire _04326_;
 wire _04327_;
 wire _04328_;
 wire _04329_;
 wire _04330_;
 wire _04331_;
 wire _04332_;
 wire _04333_;
 wire _04334_;
 wire _04335_;
 wire _04336_;
 wire _04337_;
 wire _04338_;
 wire _04339_;
 wire _04340_;
 wire _04341_;
 wire _04342_;
 wire _04343_;
 wire _04344_;
 wire _04345_;
 wire _04346_;
 wire _04347_;
 wire _04348_;
 wire _04349_;
 wire _04350_;
 wire _04351_;
 wire _04352_;
 wire _04353_;
 wire _04354_;
 wire _04355_;
 wire _04356_;
 wire _04357_;
 wire _04358_;
 wire _04359_;
 wire _04360_;
 wire _04361_;
 wire _04362_;
 wire _04363_;
 wire _04364_;
 wire _04365_;
 wire _04366_;
 wire _04367_;
 wire _04368_;
 wire _04369_;
 wire _04370_;
 wire _04371_;
 wire _04372_;
 wire _04373_;
 wire _04374_;
 wire _04375_;
 wire _04376_;
 wire _04377_;
 wire _04378_;
 wire _04379_;
 wire _04380_;
 wire _04381_;
 wire _04382_;
 wire _04383_;
 wire _04384_;
 wire _04385_;
 wire _04386_;
 wire _04387_;
 wire _04388_;
 wire _04389_;
 wire _04390_;
 wire _04391_;
 wire _04392_;
 wire _04393_;
 wire _04394_;
 wire _04395_;
 wire _04396_;
 wire _04397_;
 wire _04398_;
 wire _04399_;
 wire _04400_;
 wire _04401_;
 wire _04402_;
 wire _04403_;
 wire _04404_;
 wire _04405_;
 wire _04406_;
 wire _04407_;
 wire _04408_;
 wire _04409_;
 wire _04410_;
 wire _04411_;
 wire _04412_;
 wire _04413_;
 wire _04414_;
 wire _04415_;
 wire _04416_;
 wire _04417_;
 wire _04418_;
 wire _04419_;
 wire _04420_;
 wire _04421_;
 wire _04422_;
 wire _04423_;
 wire _04424_;
 wire _04425_;
 wire _04426_;
 wire _04427_;
 wire _04428_;
 wire _04429_;
 wire _04430_;
 wire _04431_;
 wire _04432_;
 wire _04433_;
 wire _04434_;
 wire _04435_;
 wire _04436_;
 wire _04437_;
 wire _04438_;
 wire _04439_;
 wire _04440_;
 wire _04441_;
 wire _04442_;
 wire _04443_;
 wire _04444_;
 wire _04445_;
 wire _04446_;
 wire _04447_;
 wire _04448_;
 wire _04449_;
 wire _04450_;
 wire _04451_;
 wire _04452_;
 wire _04453_;
 wire _04454_;
 wire _04455_;
 wire _04456_;
 wire _04457_;
 wire _04458_;
 wire _04459_;
 wire _04460_;
 wire _04461_;
 wire _04462_;
 wire _04463_;
 wire _04464_;
 wire _04465_;
 wire _04466_;
 wire _04467_;
 wire _04468_;
 wire _04469_;
 wire _04470_;
 wire _04471_;
 wire _04472_;
 wire _04473_;
 wire _04474_;
 wire _04475_;
 wire _04476_;
 wire _04477_;
 wire _04478_;
 wire _04479_;
 wire _04480_;
 wire _04481_;
 wire _04482_;
 wire _04483_;
 wire _04484_;
 wire _04485_;
 wire _04486_;
 wire _04487_;
 wire _04488_;
 wire _04489_;
 wire _04490_;
 wire _04491_;
 wire _04492_;
 wire _04493_;
 wire _04494_;
 wire _04495_;
 wire _04496_;
 wire _04497_;
 wire _04498_;
 wire _04499_;
 wire _04500_;
 wire _04501_;
 wire _04502_;
 wire _04503_;
 wire _04504_;
 wire _04505_;
 wire _04506_;
 wire _04507_;
 wire _04508_;
 wire _04509_;
 wire _04510_;
 wire _04511_;
 wire _04512_;
 wire _04513_;
 wire _04514_;
 wire _04515_;
 wire _04516_;
 wire _04517_;
 wire _04518_;
 wire _04519_;
 wire _04520_;
 wire _04521_;
 wire _04522_;
 wire _04523_;
 wire _04524_;
 wire _04525_;
 wire _04526_;
 wire _04527_;
 wire _04528_;
 wire _04529_;
 wire _04530_;
 wire _04531_;
 wire _04532_;
 wire _04533_;
 wire _04534_;
 wire _04535_;
 wire _04536_;
 wire _04537_;
 wire _04538_;
 wire _04539_;
 wire _04540_;
 wire _04541_;
 wire _04542_;
 wire _04543_;
 wire _04544_;
 wire _04545_;
 wire _04546_;
 wire _04547_;
 wire _04548_;
 wire _04549_;
 wire _04550_;
 wire _04551_;
 wire _04552_;
 wire _04553_;
 wire _04554_;
 wire _04555_;
 wire _04556_;
 wire _04557_;
 wire _04558_;
 wire _04559_;
 wire _04560_;
 wire _04561_;
 wire _04562_;
 wire _04563_;
 wire _04564_;
 wire _04565_;
 wire _04566_;
 wire _04567_;
 wire _04568_;
 wire _04569_;
 wire _04570_;
 wire _04571_;
 wire _04572_;
 wire _04573_;
 wire _04574_;
 wire _04575_;
 wire _04576_;
 wire _04577_;
 wire _04578_;
 wire _04579_;
 wire _04580_;
 wire _04581_;
 wire _04582_;
 wire _04583_;
 wire _04584_;
 wire _04585_;
 wire _04586_;
 wire _04587_;
 wire _04588_;
 wire _04589_;
 wire _04590_;
 wire _04591_;
 wire _04592_;
 wire _04593_;
 wire _04594_;
 wire _04595_;
 wire _04596_;
 wire _04597_;
 wire _04598_;
 wire _04599_;
 wire _04600_;
 wire _04601_;
 wire _04602_;
 wire _04603_;
 wire _04604_;
 wire _04605_;
 wire _04606_;
 wire _04607_;
 wire _04608_;
 wire _04609_;
 wire _04610_;
 wire _04611_;
 wire _04612_;
 wire _04613_;
 wire _04614_;
 wire _04615_;
 wire _04616_;
 wire _04617_;
 wire _04618_;
 wire _04619_;
 wire _04620_;
 wire _04621_;
 wire _04622_;
 wire _04623_;
 wire _04624_;
 wire _04625_;
 wire _04626_;
 wire _04627_;
 wire _04628_;
 wire _04629_;
 wire _04630_;
 wire _04631_;
 wire _04632_;
 wire _04633_;
 wire _04634_;
 wire _04635_;
 wire _04636_;
 wire _04637_;
 wire _04638_;
 wire _04639_;
 wire _04640_;
 wire _04641_;
 wire _04642_;
 wire _04643_;
 wire _04644_;
 wire _04645_;
 wire _04646_;
 wire _04647_;
 wire _04648_;
 wire _04649_;
 wire _04650_;
 wire _04651_;
 wire _04652_;
 wire _04653_;
 wire _04654_;
 wire _04655_;
 wire _04656_;
 wire _04657_;
 wire _04658_;
 wire _04659_;
 wire _04660_;
 wire _04661_;
 wire _04662_;
 wire _04663_;
 wire _04664_;
 wire _04665_;
 wire _04666_;
 wire _04667_;
 wire _04668_;
 wire _04669_;
 wire _04670_;
 wire _04671_;
 wire _04672_;
 wire _04673_;
 wire _04674_;
 wire _04675_;
 wire _04676_;
 wire _04677_;
 wire _04678_;
 wire _04679_;
 wire _04680_;
 wire _04681_;
 wire _04682_;
 wire _04683_;
 wire _04684_;
 wire _04685_;
 wire _04686_;
 wire _04687_;
 wire _04688_;
 wire _04689_;
 wire _04690_;
 wire _04691_;
 wire _04692_;
 wire _04693_;
 wire _04694_;
 wire _04695_;
 wire _04696_;
 wire _04697_;
 wire _04698_;
 wire _04699_;
 wire _04700_;
 wire _04701_;
 wire _04702_;
 wire _04703_;
 wire _04704_;
 wire _04705_;
 wire _04706_;
 wire _04707_;
 wire _04708_;
 wire _04709_;
 wire _04710_;
 wire _04711_;
 wire _04712_;
 wire _04713_;
 wire _04714_;
 wire _04715_;
 wire _04716_;
 wire _04717_;
 wire _04718_;
 wire _04719_;
 wire _04720_;
 wire _04721_;
 wire _04722_;
 wire _04723_;
 wire _04724_;
 wire _04725_;
 wire _04726_;
 wire _04727_;
 wire _04728_;
 wire _04729_;
 wire _04730_;
 wire _04731_;
 wire _04732_;
 wire _04733_;
 wire _04734_;
 wire _04735_;
 wire _04736_;
 wire _04737_;
 wire _04738_;
 wire _04739_;
 wire _04740_;
 wire _04741_;
 wire _04742_;
 wire _04743_;
 wire _04744_;
 wire _04745_;
 wire _04746_;
 wire _04747_;
 wire _04748_;
 wire _04749_;
 wire _04750_;
 wire _04751_;
 wire _04752_;
 wire _04753_;
 wire _04754_;
 wire _04755_;
 wire _04756_;
 wire _04757_;
 wire _04758_;
 wire _04759_;
 wire _04760_;
 wire _04761_;
 wire _04762_;
 wire _04763_;
 wire _04764_;
 wire _04765_;
 wire _04766_;
 wire _04767_;
 wire _04768_;
 wire _04769_;
 wire _04770_;
 wire _04771_;
 wire _04772_;
 wire _04773_;
 wire _04774_;
 wire _04775_;
 wire _04776_;
 wire _04777_;
 wire _04778_;
 wire _04779_;
 wire _04780_;
 wire _04781_;
 wire _04782_;
 wire _04783_;
 wire _04784_;
 wire _04785_;
 wire _04786_;
 wire _04787_;
 wire _04788_;
 wire _04789_;
 wire _04790_;
 wire _04791_;
 wire _04792_;
 wire _04793_;
 wire _04794_;
 wire _04795_;
 wire _04796_;
 wire _04797_;
 wire _04798_;
 wire _04799_;
 wire _04800_;
 wire _04801_;
 wire _04802_;
 wire _04803_;
 wire _04804_;
 wire _04805_;
 wire _04806_;
 wire _04807_;
 wire _04808_;
 wire _04809_;
 wire _04810_;
 wire _04811_;
 wire _04812_;
 wire _04813_;
 wire _04814_;
 wire _04815_;
 wire _04816_;
 wire _04817_;
 wire _04818_;
 wire _04819_;
 wire _04820_;
 wire _04821_;
 wire _04822_;
 wire _04823_;
 wire _04824_;
 wire _04825_;
 wire _04826_;
 wire _04827_;
 wire _04828_;
 wire _04829_;
 wire _04830_;
 wire _04831_;
 wire _04832_;
 wire _04833_;
 wire _04834_;
 wire _04835_;
 wire _04836_;
 wire _04837_;
 wire _04838_;
 wire _04839_;
 wire _04840_;
 wire _04841_;
 wire _04842_;
 wire _04843_;
 wire _04844_;
 wire _04845_;
 wire _04846_;
 wire _04847_;
 wire _04848_;
 wire _04849_;
 wire _04850_;
 wire _04851_;
 wire _04852_;
 wire _04853_;
 wire _04854_;
 wire _04855_;
 wire _04856_;
 wire _04857_;
 wire _04858_;
 wire _04859_;
 wire _04860_;
 wire _04861_;
 wire _04862_;
 wire _04863_;
 wire _04864_;
 wire _04865_;
 wire _04866_;
 wire _04867_;
 wire _04868_;
 wire _04869_;
 wire _04870_;
 wire _04871_;
 wire _04872_;
 wire _04873_;
 wire _04874_;
 wire _04875_;
 wire _04876_;
 wire _04877_;
 wire _04878_;
 wire _04879_;
 wire _04880_;
 wire _04881_;
 wire _04882_;
 wire _04883_;
 wire _04884_;
 wire _04885_;
 wire _04886_;
 wire _04887_;
 wire _04888_;
 wire _04889_;
 wire _04890_;
 wire _04891_;
 wire _04892_;
 wire _04893_;
 wire _04894_;
 wire _04895_;
 wire _04896_;
 wire _04897_;
 wire _04898_;
 wire _04899_;
 wire _04900_;
 wire _04901_;
 wire _04902_;
 wire _04903_;
 wire _04904_;
 wire _04905_;
 wire _04906_;
 wire _04907_;
 wire _04908_;
 wire _04909_;
 wire _04910_;
 wire _04911_;
 wire _04912_;
 wire _04913_;
 wire _04914_;
 wire _04915_;
 wire _04916_;
 wire _04917_;
 wire _04918_;
 wire _04919_;
 wire _04920_;
 wire _04921_;
 wire _04922_;
 wire _04923_;
 wire _04924_;
 wire _04925_;
 wire _04926_;
 wire _04927_;
 wire _04928_;
 wire _04929_;
 wire _04930_;
 wire _04931_;
 wire _04932_;
 wire _04933_;
 wire _04934_;
 wire _04935_;
 wire _04936_;
 wire _04937_;
 wire _04938_;
 wire _04939_;
 wire _04940_;
 wire _04941_;
 wire _04942_;
 wire _04943_;
 wire _04944_;
 wire _04945_;
 wire _04946_;
 wire _04947_;
 wire _04948_;
 wire _04949_;
 wire _04950_;
 wire _04951_;
 wire _04952_;
 wire _04953_;
 wire _04954_;
 wire _04955_;
 wire _04956_;
 wire _04957_;
 wire _04958_;
 wire _04959_;
 wire _04960_;
 wire _04961_;
 wire _04962_;
 wire _04963_;
 wire _04964_;
 wire _04965_;
 wire _04966_;
 wire _04967_;
 wire _04968_;
 wire _04969_;
 wire _04970_;
 wire _04971_;
 wire _04972_;
 wire _04973_;
 wire _04974_;
 wire _04975_;
 wire _04976_;
 wire _04977_;
 wire _04978_;
 wire _04979_;
 wire _04980_;
 wire _04981_;
 wire _04982_;
 wire _04983_;
 wire _04984_;
 wire _04985_;
 wire _04986_;
 wire _04987_;
 wire _04988_;
 wire _04989_;
 wire _04990_;
 wire _04991_;
 wire _04992_;
 wire _04993_;
 wire _04994_;
 wire _04995_;
 wire _04996_;
 wire _04997_;
 wire _04998_;
 wire _04999_;
 wire _05000_;
 wire _05001_;
 wire _05002_;
 wire _05003_;
 wire _05004_;
 wire _05005_;
 wire _05006_;
 wire _05007_;
 wire _05008_;
 wire _05009_;
 wire _05010_;
 wire _05011_;
 wire _05012_;
 wire _05013_;
 wire _05014_;
 wire _05015_;
 wire _05016_;
 wire _05017_;
 wire _05018_;
 wire _05019_;
 wire _05020_;
 wire _05021_;
 wire _05022_;
 wire _05023_;
 wire _05024_;
 wire _05025_;
 wire _05026_;
 wire _05027_;
 wire _05028_;
 wire _05029_;
 wire _05030_;
 wire _05031_;
 wire _05032_;
 wire _05033_;
 wire _05034_;
 wire _05035_;
 wire _05036_;
 wire _05037_;
 wire _05038_;
 wire _05039_;
 wire _05040_;
 wire _05041_;
 wire _05042_;
 wire _05043_;
 wire _05044_;
 wire _05045_;
 wire _05046_;
 wire _05047_;
 wire _05048_;
 wire _05049_;
 wire _05050_;
 wire _05051_;
 wire _05052_;
 wire _05053_;
 wire _05054_;
 wire _05055_;
 wire _05056_;
 wire _05057_;
 wire _05058_;
 wire _05059_;
 wire _05060_;
 wire _05061_;
 wire _05062_;
 wire _05063_;
 wire _05064_;
 wire _05065_;
 wire _05066_;
 wire _05067_;
 wire _05068_;
 wire _05069_;
 wire _05070_;
 wire _05071_;
 wire _05072_;
 wire _05073_;
 wire _05074_;
 wire _05075_;
 wire _05076_;
 wire _05077_;
 wire _05078_;
 wire _05079_;
 wire _05080_;
 wire _05081_;
 wire _05082_;
 wire _05083_;
 wire _05084_;
 wire _05085_;
 wire _05086_;
 wire _05087_;
 wire _05088_;
 wire _05089_;
 wire _05090_;
 wire _05091_;
 wire _05092_;
 wire _05093_;
 wire _05094_;
 wire _05095_;
 wire _05096_;
 wire _05097_;
 wire _05098_;
 wire _05099_;
 wire _05100_;
 wire _05101_;
 wire _05102_;
 wire _05103_;
 wire _05104_;
 wire _05105_;
 wire _05106_;
 wire _05107_;
 wire _05108_;
 wire _05109_;
 wire _05110_;
 wire _05111_;
 wire _05112_;
 wire _05113_;
 wire _05114_;
 wire _05115_;
 wire _05116_;
 wire _05117_;
 wire _05118_;
 wire _05119_;
 wire _05120_;
 wire _05121_;
 wire _05122_;
 wire _05123_;
 wire _05124_;
 wire _05125_;
 wire _05126_;
 wire _05127_;
 wire _05128_;
 wire _05129_;
 wire _05130_;
 wire _05131_;
 wire _05132_;
 wire _05133_;
 wire _05134_;
 wire _05135_;
 wire _05136_;
 wire _05137_;
 wire _05138_;
 wire _05139_;
 wire _05140_;
 wire _05141_;
 wire _05142_;
 wire _05143_;
 wire _05144_;
 wire _05145_;
 wire _05146_;
 wire _05147_;
 wire _05148_;
 wire _05149_;
 wire _05150_;
 wire _05151_;
 wire _05152_;
 wire _05153_;
 wire _05154_;
 wire _05155_;
 wire _05156_;
 wire _05157_;
 wire _05158_;
 wire _05159_;
 wire _05160_;
 wire _05161_;
 wire _05162_;
 wire _05163_;
 wire _05164_;
 wire _05165_;
 wire _05166_;
 wire _05167_;
 wire _05168_;
 wire _05169_;
 wire _05170_;
 wire _05171_;
 wire _05172_;
 wire _05173_;
 wire _05174_;
 wire _05175_;
 wire _05176_;
 wire _05177_;
 wire _05178_;
 wire _05179_;
 wire _05180_;
 wire _05181_;
 wire _05182_;
 wire _05183_;
 wire _05184_;
 wire _05185_;
 wire _05186_;
 wire _05187_;
 wire _05188_;
 wire _05189_;
 wire _05190_;
 wire _05191_;
 wire _05192_;
 wire _05193_;
 wire _05194_;
 wire _05195_;
 wire _05196_;
 wire _05197_;
 wire _05198_;
 wire _05199_;
 wire _05200_;
 wire _05201_;
 wire _05202_;
 wire _05203_;
 wire _05204_;
 wire _05205_;
 wire _05206_;
 wire _05207_;
 wire _05208_;
 wire _05209_;
 wire _05210_;
 wire _05211_;
 wire _05212_;
 wire _05213_;
 wire _05214_;
 wire _05215_;
 wire _05216_;
 wire _05217_;
 wire _05218_;
 wire _05219_;
 wire _05220_;
 wire _05221_;
 wire _05222_;
 wire _05223_;
 wire _05224_;
 wire _05225_;
 wire _05226_;
 wire _05227_;
 wire _05228_;
 wire _05229_;
 wire _05230_;
 wire _05231_;
 wire _05232_;
 wire _05233_;
 wire _05234_;
 wire _05235_;
 wire _05236_;
 wire _05237_;
 wire _05238_;
 wire _05239_;
 wire _05240_;
 wire _05241_;
 wire _05242_;
 wire _05243_;
 wire _05244_;
 wire _05245_;
 wire _05246_;
 wire _05247_;
 wire _05248_;
 wire _05249_;
 wire _05250_;
 wire _05251_;
 wire _05252_;
 wire _05253_;
 wire _05254_;
 wire _05255_;
 wire _05256_;
 wire _05257_;
 wire _05258_;
 wire _05259_;
 wire _05260_;
 wire _05261_;
 wire _05262_;
 wire _05263_;
 wire _05264_;
 wire _05265_;
 wire _05266_;
 wire _05267_;
 wire _05268_;
 wire _05269_;
 wire _05270_;
 wire _05271_;
 wire _05272_;
 wire _05273_;
 wire _05274_;
 wire _05275_;
 wire _05276_;
 wire _05277_;
 wire _05278_;
 wire _05279_;
 wire _05280_;
 wire _05281_;
 wire _05282_;
 wire _05283_;
 wire _05284_;
 wire _05285_;
 wire _05286_;
 wire _05287_;
 wire _05288_;
 wire _05289_;
 wire _05290_;
 wire _05291_;
 wire _05292_;
 wire _05293_;
 wire _05294_;
 wire _05295_;
 wire _05296_;
 wire _05297_;
 wire _05298_;
 wire _05299_;
 wire _05300_;
 wire _05301_;
 wire _05302_;
 wire _05303_;
 wire _05304_;
 wire _05305_;
 wire _05306_;
 wire _05307_;
 wire _05308_;
 wire _05309_;
 wire _05310_;
 wire _05311_;
 wire _05312_;
 wire _05313_;
 wire _05314_;
 wire _05315_;
 wire _05316_;
 wire _05317_;
 wire _05318_;
 wire _05319_;
 wire _05320_;
 wire _05321_;
 wire _05322_;
 wire _05323_;
 wire _05324_;
 wire _05325_;
 wire _05326_;
 wire _05327_;
 wire _05328_;
 wire _05329_;
 wire _05330_;
 wire _05331_;
 wire _05332_;
 wire _05333_;
 wire _05334_;
 wire _05335_;
 wire _05336_;
 wire _05337_;
 wire _05338_;
 wire _05339_;
 wire _05340_;
 wire _05341_;
 wire _05342_;
 wire _05343_;
 wire _05344_;
 wire _05345_;
 wire _05346_;
 wire _05347_;
 wire _05348_;
 wire _05349_;
 wire _05350_;
 wire _05351_;
 wire _05352_;
 wire _05353_;
 wire _05354_;
 wire _05355_;
 wire _05356_;
 wire _05357_;
 wire _05358_;
 wire _05359_;
 wire _05360_;
 wire _05361_;
 wire _05362_;
 wire _05363_;
 wire _05364_;
 wire _05365_;
 wire _05366_;
 wire _05367_;
 wire _05368_;
 wire _05369_;
 wire _05370_;
 wire _05371_;
 wire _05372_;
 wire _05373_;
 wire _05374_;
 wire _05375_;
 wire _05376_;
 wire _05377_;
 wire _05378_;
 wire _05379_;
 wire _05380_;
 wire _05381_;
 wire _05382_;
 wire _05383_;
 wire _05384_;
 wire _05385_;
 wire _05386_;
 wire _05387_;
 wire _05388_;
 wire _05389_;
 wire _05390_;
 wire _05391_;
 wire _05392_;
 wire _05393_;
 wire _05394_;
 wire _05395_;
 wire _05396_;
 wire _05397_;
 wire _05398_;
 wire _05399_;
 wire _05400_;
 wire _05401_;
 wire _05402_;
 wire _05403_;
 wire _05404_;
 wire _05405_;
 wire _05406_;
 wire _05407_;
 wire _05408_;
 wire _05409_;
 wire _05410_;
 wire _05411_;
 wire _05412_;
 wire _05413_;
 wire _05414_;
 wire _05415_;
 wire _05416_;
 wire _05417_;
 wire _05418_;
 wire _05419_;
 wire _05420_;
 wire _05421_;
 wire _05422_;
 wire _05423_;
 wire _05424_;
 wire _05425_;
 wire _05426_;
 wire _05427_;
 wire _05428_;
 wire _05429_;
 wire _05430_;
 wire _05431_;
 wire _05432_;
 wire _05433_;
 wire _05434_;
 wire _05435_;
 wire _05436_;
 wire _05437_;
 wire _05438_;
 wire _05439_;
 wire _05440_;
 wire _05441_;
 wire _05442_;
 wire _05443_;
 wire _05444_;
 wire _05445_;
 wire _05446_;
 wire _05447_;
 wire _05448_;
 wire _05449_;
 wire _05450_;
 wire _05451_;
 wire _05452_;
 wire _05453_;
 wire _05454_;
 wire _05455_;
 wire _05456_;
 wire _05457_;
 wire _05458_;
 wire _05459_;
 wire _05460_;
 wire _05461_;
 wire net92;
 wire net102;
 wire net103;
 wire net93;
 wire net104;
 wire net105;
 wire net225;
 wire net106;
 wire net107;
 wire net108;
 wire net94;
 wire net226;
 wire net227;
 wire net228;
 wire clknet_leaf_0_wb_clk_i;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net113;
 wire net114;
 wire net121;
 wire net115;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net130;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net131;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net132;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net133;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net134;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire \soc.boot_loading_offset[0] ;
 wire \soc.boot_loading_offset[1] ;
 wire \soc.boot_loading_offset[2] ;
 wire \soc.boot_loading_offset[3] ;
 wire \soc.boot_loading_offset[4] ;
 wire \soc.cpu.ALU.f ;
 wire \soc.cpu.ALU.no ;
 wire \soc.cpu.ALU.nx ;
 wire \soc.cpu.ALU.ny ;
 wire \soc.cpu.ALU.x[0] ;
 wire \soc.cpu.ALU.x[10] ;
 wire \soc.cpu.ALU.x[11] ;
 wire \soc.cpu.ALU.x[12] ;
 wire \soc.cpu.ALU.x[13] ;
 wire \soc.cpu.ALU.x[14] ;
 wire \soc.cpu.ALU.x[15] ;
 wire \soc.cpu.ALU.x[1] ;
 wire \soc.cpu.ALU.x[2] ;
 wire \soc.cpu.ALU.x[3] ;
 wire \soc.cpu.ALU.x[4] ;
 wire \soc.cpu.ALU.x[5] ;
 wire \soc.cpu.ALU.x[6] ;
 wire \soc.cpu.ALU.x[7] ;
 wire \soc.cpu.ALU.x[8] ;
 wire \soc.cpu.ALU.x[9] ;
 wire \soc.cpu.ALU.zx ;
 wire \soc.cpu.ALU.zy ;
 wire \soc.cpu.AReg.clk ;
 wire \soc.cpu.AReg.data[0] ;
 wire \soc.cpu.AReg.data[10] ;
 wire \soc.cpu.AReg.data[11] ;
 wire \soc.cpu.AReg.data[12] ;
 wire \soc.cpu.AReg.data[13] ;
 wire \soc.cpu.AReg.data[14] ;
 wire \soc.cpu.AReg.data[15] ;
 wire \soc.cpu.AReg.data[1] ;
 wire \soc.cpu.AReg.data[2] ;
 wire \soc.cpu.AReg.data[3] ;
 wire \soc.cpu.AReg.data[4] ;
 wire \soc.cpu.AReg.data[5] ;
 wire \soc.cpu.AReg.data[6] ;
 wire \soc.cpu.AReg.data[7] ;
 wire \soc.cpu.AReg.data[8] ;
 wire \soc.cpu.AReg.data[9] ;
 wire \soc.cpu.DMuxJMP.sel[0] ;
 wire \soc.cpu.DMuxJMP.sel[1] ;
 wire \soc.cpu.DMuxJMP.sel[2] ;
 wire \soc.cpu.PC.REG.data[0] ;
 wire \soc.cpu.PC.REG.data[10] ;
 wire \soc.cpu.PC.REG.data[11] ;
 wire \soc.cpu.PC.REG.data[12] ;
 wire \soc.cpu.PC.REG.data[13] ;
 wire \soc.cpu.PC.REG.data[14] ;
 wire \soc.cpu.PC.REG.data[1] ;
 wire \soc.cpu.PC.REG.data[2] ;
 wire \soc.cpu.PC.REG.data[3] ;
 wire \soc.cpu.PC.REG.data[4] ;
 wire \soc.cpu.PC.REG.data[5] ;
 wire \soc.cpu.PC.REG.data[6] ;
 wire \soc.cpu.PC.REG.data[7] ;
 wire \soc.cpu.PC.REG.data[8] ;
 wire \soc.cpu.PC.REG.data[9] ;
 wire \soc.cpu.PC.in[0] ;
 wire \soc.cpu.PC.in[10] ;
 wire \soc.cpu.PC.in[11] ;
 wire \soc.cpu.PC.in[12] ;
 wire \soc.cpu.PC.in[13] ;
 wire \soc.cpu.PC.in[14] ;
 wire \soc.cpu.PC.in[1] ;
 wire \soc.cpu.PC.in[2] ;
 wire \soc.cpu.PC.in[3] ;
 wire \soc.cpu.PC.in[4] ;
 wire \soc.cpu.PC.in[5] ;
 wire \soc.cpu.PC.in[6] ;
 wire \soc.cpu.PC.in[7] ;
 wire \soc.cpu.PC.in[8] ;
 wire \soc.cpu.PC.in[9] ;
 wire \soc.cpu.instruction[12] ;
 wire \soc.cpu.instruction[13] ;
 wire \soc.cpu.instruction[14] ;
 wire \soc.cpu.instruction[15] ;
 wire \soc.cpu.instruction[3] ;
 wire \soc.cpu.instruction[4] ;
 wire \soc.cpu.instruction[5] ;
 wire \soc.display_clks_before_active[0] ;
 wire \soc.gpio_i_stored[0] ;
 wire \soc.gpio_i_stored[1] ;
 wire \soc.gpio_i_stored[2] ;
 wire \soc.gpio_i_stored[3] ;
 wire \soc.hack_clk_strobe ;
 wire \soc.hack_clock_0.counter[0] ;
 wire \soc.hack_clock_0.counter[1] ;
 wire \soc.hack_clock_0.counter[2] ;
 wire \soc.hack_clock_0.counter[3] ;
 wire \soc.hack_clock_0.counter[4] ;
 wire \soc.hack_clock_0.counter[5] ;
 wire \soc.hack_clock_0.counter[6] ;
 wire \soc.hack_rom_request ;
 wire \soc.hack_wait_clocks[0] ;
 wire \soc.hack_wait_clocks[1] ;
 wire \soc.ram_data_out[0] ;
 wire \soc.ram_data_out[10] ;
 wire \soc.ram_data_out[11] ;
 wire \soc.ram_data_out[12] ;
 wire \soc.ram_data_out[13] ;
 wire \soc.ram_data_out[14] ;
 wire \soc.ram_data_out[15] ;
 wire \soc.ram_data_out[1] ;
 wire \soc.ram_data_out[2] ;
 wire \soc.ram_data_out[3] ;
 wire \soc.ram_data_out[4] ;
 wire \soc.ram_data_out[5] ;
 wire \soc.ram_data_out[6] ;
 wire \soc.ram_data_out[7] ;
 wire \soc.ram_data_out[8] ;
 wire \soc.ram_data_out[9] ;
 wire \soc.ram_encoder_0.address[0] ;
 wire \soc.ram_encoder_0.address[10] ;
 wire \soc.ram_encoder_0.address[11] ;
 wire \soc.ram_encoder_0.address[12] ;
 wire \soc.ram_encoder_0.address[13] ;
 wire \soc.ram_encoder_0.address[14] ;
 wire \soc.ram_encoder_0.address[1] ;
 wire \soc.ram_encoder_0.address[2] ;
 wire \soc.ram_encoder_0.address[3] ;
 wire \soc.ram_encoder_0.address[4] ;
 wire \soc.ram_encoder_0.address[5] ;
 wire \soc.ram_encoder_0.address[6] ;
 wire \soc.ram_encoder_0.address[7] ;
 wire \soc.ram_encoder_0.address[8] ;
 wire \soc.ram_encoder_0.address[9] ;
 wire \soc.ram_encoder_0.current_state[0] ;
 wire \soc.ram_encoder_0.current_state[1] ;
 wire \soc.ram_encoder_0.current_state[2] ;
 wire \soc.ram_encoder_0.data_out[0] ;
 wire \soc.ram_encoder_0.data_out[10] ;
 wire \soc.ram_encoder_0.data_out[11] ;
 wire \soc.ram_encoder_0.data_out[12] ;
 wire \soc.ram_encoder_0.data_out[13] ;
 wire \soc.ram_encoder_0.data_out[14] ;
 wire \soc.ram_encoder_0.data_out[15] ;
 wire \soc.ram_encoder_0.data_out[1] ;
 wire \soc.ram_encoder_0.data_out[2] ;
 wire \soc.ram_encoder_0.data_out[3] ;
 wire \soc.ram_encoder_0.data_out[4] ;
 wire \soc.ram_encoder_0.data_out[5] ;
 wire \soc.ram_encoder_0.data_out[6] ;
 wire \soc.ram_encoder_0.data_out[7] ;
 wire \soc.ram_encoder_0.data_out[8] ;
 wire \soc.ram_encoder_0.data_out[9] ;
 wire \soc.ram_encoder_0.initialized ;
 wire \soc.ram_encoder_0.initializing_step[0] ;
 wire \soc.ram_encoder_0.initializing_step[1] ;
 wire \soc.ram_encoder_0.initializing_step[2] ;
 wire \soc.ram_encoder_0.initializing_step[3] ;
 wire \soc.ram_encoder_0.initializing_step[4] ;
 wire \soc.ram_encoder_0.input_bits_left[2] ;
 wire \soc.ram_encoder_0.input_bits_left[3] ;
 wire \soc.ram_encoder_0.input_bits_left[4] ;
 wire \soc.ram_encoder_0.input_buffer[0] ;
 wire \soc.ram_encoder_0.input_buffer[10] ;
 wire \soc.ram_encoder_0.input_buffer[11] ;
 wire \soc.ram_encoder_0.input_buffer[1] ;
 wire \soc.ram_encoder_0.input_buffer[2] ;
 wire \soc.ram_encoder_0.input_buffer[3] ;
 wire \soc.ram_encoder_0.input_buffer[4] ;
 wire \soc.ram_encoder_0.input_buffer[5] ;
 wire \soc.ram_encoder_0.input_buffer[6] ;
 wire \soc.ram_encoder_0.input_buffer[7] ;
 wire \soc.ram_encoder_0.input_buffer[8] ;
 wire \soc.ram_encoder_0.input_buffer[9] ;
 wire \soc.ram_encoder_0.output_bits_left[2] ;
 wire \soc.ram_encoder_0.output_bits_left[3] ;
 wire \soc.ram_encoder_0.output_bits_left[4] ;
 wire \soc.ram_encoder_0.output_buffer[10] ;
 wire \soc.ram_encoder_0.output_buffer[11] ;
 wire \soc.ram_encoder_0.output_buffer[12] ;
 wire \soc.ram_encoder_0.output_buffer[13] ;
 wire \soc.ram_encoder_0.output_buffer[14] ;
 wire \soc.ram_encoder_0.output_buffer[15] ;
 wire \soc.ram_encoder_0.output_buffer[16] ;
 wire \soc.ram_encoder_0.output_buffer[17] ;
 wire \soc.ram_encoder_0.output_buffer[18] ;
 wire \soc.ram_encoder_0.output_buffer[19] ;
 wire \soc.ram_encoder_0.output_buffer[1] ;
 wire \soc.ram_encoder_0.output_buffer[2] ;
 wire \soc.ram_encoder_0.output_buffer[3] ;
 wire \soc.ram_encoder_0.output_buffer[4] ;
 wire \soc.ram_encoder_0.output_buffer[5] ;
 wire \soc.ram_encoder_0.output_buffer[6] ;
 wire \soc.ram_encoder_0.output_buffer[7] ;
 wire \soc.ram_encoder_0.output_buffer[8] ;
 wire \soc.ram_encoder_0.output_buffer[9] ;
 wire \soc.ram_encoder_0.request_address[0] ;
 wire \soc.ram_encoder_0.request_address[10] ;
 wire \soc.ram_encoder_0.request_address[11] ;
 wire \soc.ram_encoder_0.request_address[12] ;
 wire \soc.ram_encoder_0.request_address[13] ;
 wire \soc.ram_encoder_0.request_address[14] ;
 wire \soc.ram_encoder_0.request_address[1] ;
 wire \soc.ram_encoder_0.request_address[2] ;
 wire \soc.ram_encoder_0.request_address[3] ;
 wire \soc.ram_encoder_0.request_address[4] ;
 wire \soc.ram_encoder_0.request_address[5] ;
 wire \soc.ram_encoder_0.request_address[6] ;
 wire \soc.ram_encoder_0.request_address[7] ;
 wire \soc.ram_encoder_0.request_address[8] ;
 wire \soc.ram_encoder_0.request_address[9] ;
 wire \soc.ram_encoder_0.request_data_out[0] ;
 wire \soc.ram_encoder_0.request_data_out[10] ;
 wire \soc.ram_encoder_0.request_data_out[11] ;
 wire \soc.ram_encoder_0.request_data_out[12] ;
 wire \soc.ram_encoder_0.request_data_out[13] ;
 wire \soc.ram_encoder_0.request_data_out[14] ;
 wire \soc.ram_encoder_0.request_data_out[15] ;
 wire \soc.ram_encoder_0.request_data_out[1] ;
 wire \soc.ram_encoder_0.request_data_out[2] ;
 wire \soc.ram_encoder_0.request_data_out[3] ;
 wire \soc.ram_encoder_0.request_data_out[4] ;
 wire \soc.ram_encoder_0.request_data_out[5] ;
 wire \soc.ram_encoder_0.request_data_out[6] ;
 wire \soc.ram_encoder_0.request_data_out[7] ;
 wire \soc.ram_encoder_0.request_data_out[8] ;
 wire \soc.ram_encoder_0.request_data_out[9] ;
 wire \soc.ram_encoder_0.request_write ;
 wire \soc.ram_encoder_0.sram_sio_oe ;
 wire \soc.ram_encoder_0.toggled_sram_sck ;
 wire \soc.ram_step1_write_request ;
 wire \soc.ram_step2_read_request ;
 wire \soc.rom_encoder_0.current_state[0] ;
 wire \soc.rom_encoder_0.current_state[1] ;
 wire \soc.rom_encoder_0.current_state[2] ;
 wire \soc.rom_encoder_0.data_out[0] ;
 wire \soc.rom_encoder_0.data_out[10] ;
 wire \soc.rom_encoder_0.data_out[11] ;
 wire \soc.rom_encoder_0.data_out[12] ;
 wire \soc.rom_encoder_0.data_out[13] ;
 wire \soc.rom_encoder_0.data_out[14] ;
 wire \soc.rom_encoder_0.data_out[15] ;
 wire \soc.rom_encoder_0.data_out[1] ;
 wire \soc.rom_encoder_0.data_out[2] ;
 wire \soc.rom_encoder_0.data_out[3] ;
 wire \soc.rom_encoder_0.data_out[4] ;
 wire \soc.rom_encoder_0.data_out[5] ;
 wire \soc.rom_encoder_0.data_out[6] ;
 wire \soc.rom_encoder_0.data_out[7] ;
 wire \soc.rom_encoder_0.data_out[8] ;
 wire \soc.rom_encoder_0.data_out[9] ;
 wire \soc.rom_encoder_0.initialized ;
 wire \soc.rom_encoder_0.initializing_step[0] ;
 wire \soc.rom_encoder_0.initializing_step[1] ;
 wire \soc.rom_encoder_0.initializing_step[2] ;
 wire \soc.rom_encoder_0.initializing_step[3] ;
 wire \soc.rom_encoder_0.initializing_step[4] ;
 wire \soc.rom_encoder_0.input_bits_left[2] ;
 wire \soc.rom_encoder_0.input_bits_left[3] ;
 wire \soc.rom_encoder_0.input_bits_left[4] ;
 wire \soc.rom_encoder_0.input_buffer[0] ;
 wire \soc.rom_encoder_0.input_buffer[10] ;
 wire \soc.rom_encoder_0.input_buffer[11] ;
 wire \soc.rom_encoder_0.input_buffer[1] ;
 wire \soc.rom_encoder_0.input_buffer[2] ;
 wire \soc.rom_encoder_0.input_buffer[3] ;
 wire \soc.rom_encoder_0.input_buffer[4] ;
 wire \soc.rom_encoder_0.input_buffer[5] ;
 wire \soc.rom_encoder_0.input_buffer[6] ;
 wire \soc.rom_encoder_0.input_buffer[7] ;
 wire \soc.rom_encoder_0.input_buffer[8] ;
 wire \soc.rom_encoder_0.input_buffer[9] ;
 wire \soc.rom_encoder_0.output_bits_left[2] ;
 wire \soc.rom_encoder_0.output_bits_left[3] ;
 wire \soc.rom_encoder_0.output_bits_left[4] ;
 wire \soc.rom_encoder_0.output_buffer[10] ;
 wire \soc.rom_encoder_0.output_buffer[11] ;
 wire \soc.rom_encoder_0.output_buffer[12] ;
 wire \soc.rom_encoder_0.output_buffer[13] ;
 wire \soc.rom_encoder_0.output_buffer[14] ;
 wire \soc.rom_encoder_0.output_buffer[15] ;
 wire \soc.rom_encoder_0.output_buffer[16] ;
 wire \soc.rom_encoder_0.output_buffer[17] ;
 wire \soc.rom_encoder_0.output_buffer[18] ;
 wire \soc.rom_encoder_0.output_buffer[19] ;
 wire \soc.rom_encoder_0.output_buffer[1] ;
 wire \soc.rom_encoder_0.output_buffer[2] ;
 wire \soc.rom_encoder_0.output_buffer[3] ;
 wire \soc.rom_encoder_0.output_buffer[4] ;
 wire \soc.rom_encoder_0.output_buffer[5] ;
 wire \soc.rom_encoder_0.output_buffer[6] ;
 wire \soc.rom_encoder_0.output_buffer[7] ;
 wire \soc.rom_encoder_0.output_buffer[8] ;
 wire \soc.rom_encoder_0.output_buffer[9] ;
 wire \soc.rom_encoder_0.request_address[0] ;
 wire \soc.rom_encoder_0.request_address[10] ;
 wire \soc.rom_encoder_0.request_address[11] ;
 wire \soc.rom_encoder_0.request_address[12] ;
 wire \soc.rom_encoder_0.request_address[13] ;
 wire \soc.rom_encoder_0.request_address[14] ;
 wire \soc.rom_encoder_0.request_address[1] ;
 wire \soc.rom_encoder_0.request_address[2] ;
 wire \soc.rom_encoder_0.request_address[3] ;
 wire \soc.rom_encoder_0.request_address[4] ;
 wire \soc.rom_encoder_0.request_address[5] ;
 wire \soc.rom_encoder_0.request_address[6] ;
 wire \soc.rom_encoder_0.request_address[7] ;
 wire \soc.rom_encoder_0.request_address[8] ;
 wire \soc.rom_encoder_0.request_address[9] ;
 wire \soc.rom_encoder_0.request_data_out[0] ;
 wire \soc.rom_encoder_0.request_data_out[10] ;
 wire \soc.rom_encoder_0.request_data_out[11] ;
 wire \soc.rom_encoder_0.request_data_out[12] ;
 wire \soc.rom_encoder_0.request_data_out[13] ;
 wire \soc.rom_encoder_0.request_data_out[14] ;
 wire \soc.rom_encoder_0.request_data_out[15] ;
 wire \soc.rom_encoder_0.request_data_out[1] ;
 wire \soc.rom_encoder_0.request_data_out[2] ;
 wire \soc.rom_encoder_0.request_data_out[3] ;
 wire \soc.rom_encoder_0.request_data_out[4] ;
 wire \soc.rom_encoder_0.request_data_out[5] ;
 wire \soc.rom_encoder_0.request_data_out[6] ;
 wire \soc.rom_encoder_0.request_data_out[7] ;
 wire \soc.rom_encoder_0.request_data_out[8] ;
 wire \soc.rom_encoder_0.request_data_out[9] ;
 wire \soc.rom_encoder_0.request_write ;
 wire \soc.rom_encoder_0.sram_sio_oe ;
 wire \soc.rom_encoder_0.toggled_sram_sck ;
 wire \soc.rom_encoder_0.write_enable ;
 wire \soc.rom_loader.current_address[0] ;
 wire \soc.rom_loader.current_address[10] ;
 wire \soc.rom_loader.current_address[11] ;
 wire \soc.rom_loader.current_address[12] ;
 wire \soc.rom_loader.current_address[13] ;
 wire \soc.rom_loader.current_address[14] ;
 wire \soc.rom_loader.current_address[1] ;
 wire \soc.rom_loader.current_address[2] ;
 wire \soc.rom_loader.current_address[3] ;
 wire \soc.rom_loader.current_address[4] ;
 wire \soc.rom_loader.current_address[5] ;
 wire \soc.rom_loader.current_address[6] ;
 wire \soc.rom_loader.current_address[7] ;
 wire \soc.rom_loader.current_address[8] ;
 wire \soc.rom_loader.current_address[9] ;
 wire \soc.rom_loader.rom_request ;
 wire \soc.rom_loader.wait_fall_clk ;
 wire \soc.rom_loader.was_loading ;
 wire \soc.rom_loader.writing ;
 wire \soc.spi_video_ram_1.buffer_index[0] ;
 wire \soc.spi_video_ram_1.buffer_index[1] ;
 wire \soc.spi_video_ram_1.buffer_index[2] ;
 wire \soc.spi_video_ram_1.buffer_index[3] ;
 wire \soc.spi_video_ram_1.buffer_index[4] ;
 wire \soc.spi_video_ram_1.buffer_index[5] ;
 wire \soc.spi_video_ram_1.current_state[0] ;
 wire \soc.spi_video_ram_1.current_state[1] ;
 wire \soc.spi_video_ram_1.current_state[2] ;
 wire \soc.spi_video_ram_1.current_state[3] ;
 wire \soc.spi_video_ram_1.current_state[4] ;
 wire \soc.spi_video_ram_1.fifo_in_address[0] ;
 wire \soc.spi_video_ram_1.fifo_in_address[10] ;
 wire \soc.spi_video_ram_1.fifo_in_address[11] ;
 wire \soc.spi_video_ram_1.fifo_in_address[12] ;
 wire \soc.spi_video_ram_1.fifo_in_address[1] ;
 wire \soc.spi_video_ram_1.fifo_in_address[2] ;
 wire \soc.spi_video_ram_1.fifo_in_address[3] ;
 wire \soc.spi_video_ram_1.fifo_in_address[4] ;
 wire \soc.spi_video_ram_1.fifo_in_address[5] ;
 wire \soc.spi_video_ram_1.fifo_in_address[6] ;
 wire \soc.spi_video_ram_1.fifo_in_address[7] ;
 wire \soc.spi_video_ram_1.fifo_in_address[8] ;
 wire \soc.spi_video_ram_1.fifo_in_address[9] ;
 wire \soc.spi_video_ram_1.fifo_in_data[0] ;
 wire \soc.spi_video_ram_1.fifo_in_data[10] ;
 wire \soc.spi_video_ram_1.fifo_in_data[11] ;
 wire \soc.spi_video_ram_1.fifo_in_data[12] ;
 wire \soc.spi_video_ram_1.fifo_in_data[13] ;
 wire \soc.spi_video_ram_1.fifo_in_data[14] ;
 wire \soc.spi_video_ram_1.fifo_in_data[15] ;
 wire \soc.spi_video_ram_1.fifo_in_data[1] ;
 wire \soc.spi_video_ram_1.fifo_in_data[2] ;
 wire \soc.spi_video_ram_1.fifo_in_data[3] ;
 wire \soc.spi_video_ram_1.fifo_in_data[4] ;
 wire \soc.spi_video_ram_1.fifo_in_data[5] ;
 wire \soc.spi_video_ram_1.fifo_in_data[6] ;
 wire \soc.spi_video_ram_1.fifo_in_data[7] ;
 wire \soc.spi_video_ram_1.fifo_in_data[8] ;
 wire \soc.spi_video_ram_1.fifo_in_data[9] ;
 wire \soc.spi_video_ram_1.fifo_read_request ;
 wire \soc.spi_video_ram_1.fifo_write_request ;
 wire \soc.spi_video_ram_1.initialized ;
 wire \soc.spi_video_ram_1.output_buffer[10] ;
 wire \soc.spi_video_ram_1.output_buffer[11] ;
 wire \soc.spi_video_ram_1.output_buffer[12] ;
 wire \soc.spi_video_ram_1.output_buffer[13] ;
 wire \soc.spi_video_ram_1.output_buffer[14] ;
 wire \soc.spi_video_ram_1.output_buffer[15] ;
 wire \soc.spi_video_ram_1.output_buffer[16] ;
 wire \soc.spi_video_ram_1.output_buffer[17] ;
 wire \soc.spi_video_ram_1.output_buffer[18] ;
 wire \soc.spi_video_ram_1.output_buffer[19] ;
 wire \soc.spi_video_ram_1.output_buffer[1] ;
 wire \soc.spi_video_ram_1.output_buffer[20] ;
 wire \soc.spi_video_ram_1.output_buffer[21] ;
 wire \soc.spi_video_ram_1.output_buffer[22] ;
 wire \soc.spi_video_ram_1.output_buffer[23] ;
 wire \soc.spi_video_ram_1.output_buffer[2] ;
 wire \soc.spi_video_ram_1.output_buffer[3] ;
 wire \soc.spi_video_ram_1.output_buffer[4] ;
 wire \soc.spi_video_ram_1.output_buffer[5] ;
 wire \soc.spi_video_ram_1.output_buffer[6] ;
 wire \soc.spi_video_ram_1.output_buffer[7] ;
 wire \soc.spi_video_ram_1.output_buffer[8] ;
 wire \soc.spi_video_ram_1.output_buffer[9] ;
 wire \soc.spi_video_ram_1.read_value[0] ;
 wire \soc.spi_video_ram_1.read_value[1] ;
 wire \soc.spi_video_ram_1.read_value[2] ;
 wire \soc.spi_video_ram_1.read_value[3] ;
 wire \soc.spi_video_ram_1.sram_sck_fall_edge ;
 wire \soc.spi_video_ram_1.sram_sck_rise_edge ;
 wire \soc.spi_video_ram_1.sram_sio_oe ;
 wire \soc.spi_video_ram_1.start_read ;
 wire \soc.spi_video_ram_1.state_counter[0] ;
 wire \soc.spi_video_ram_1.state_counter[10] ;
 wire \soc.spi_video_ram_1.state_counter[1] ;
 wire \soc.spi_video_ram_1.state_counter[2] ;
 wire \soc.spi_video_ram_1.state_counter[3] ;
 wire \soc.spi_video_ram_1.state_counter[4] ;
 wire \soc.spi_video_ram_1.state_counter[5] ;
 wire \soc.spi_video_ram_1.state_counter[6] ;
 wire \soc.spi_video_ram_1.state_counter[7] ;
 wire \soc.spi_video_ram_1.state_counter[8] ;
 wire \soc.spi_video_ram_1.state_counter[9] ;
 wire \soc.spi_video_ram_1.state_sram_clk_counter[0] ;
 wire \soc.spi_video_ram_1.state_sram_clk_counter[1] ;
 wire \soc.spi_video_ram_1.state_sram_clk_counter[2] ;
 wire \soc.spi_video_ram_1.state_sram_clk_counter[3] ;
 wire \soc.spi_video_ram_1.state_sram_clk_counter[4] ;
 wire \soc.spi_video_ram_1.state_sram_clk_counter[5] ;
 wire \soc.spi_video_ram_1.state_sram_clk_counter[6] ;
 wire \soc.spi_video_ram_1.state_sram_clk_counter[7] ;
 wire \soc.spi_video_ram_1.state_sram_clk_counter[8] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[0][0] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[0][10] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[0][11] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[0][12] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[0][13] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[0][14] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[0][15] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[0][16] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[0][17] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[0][18] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[0][19] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[0][1] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[0][20] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[0][21] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[0][22] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[0][23] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[0][24] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[0][25] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[0][26] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[0][27] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[0][28] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[0][2] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[0][3] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[0][4] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[0][5] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[0][6] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[0][7] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[0][8] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[0][9] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[10][0] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[10][10] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[10][11] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[10][12] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[10][13] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[10][14] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[10][15] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[10][16] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[10][17] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[10][18] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[10][19] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[10][1] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[10][20] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[10][21] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[10][22] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[10][23] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[10][24] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[10][25] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[10][26] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[10][27] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[10][28] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[10][2] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[10][3] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[10][4] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[10][5] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[10][6] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[10][7] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[10][8] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[10][9] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[11][0] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[11][10] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[11][11] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[11][12] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[11][13] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[11][14] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[11][15] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[11][16] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[11][17] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[11][18] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[11][19] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[11][1] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[11][20] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[11][21] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[11][22] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[11][23] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[11][24] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[11][25] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[11][26] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[11][27] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[11][28] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[11][2] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[11][3] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[11][4] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[11][5] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[11][6] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[11][7] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[11][8] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[11][9] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[12][0] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[12][10] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[12][11] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[12][12] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[12][13] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[12][14] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[12][15] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[12][16] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[12][17] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[12][18] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[12][19] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[12][1] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[12][20] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[12][21] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[12][22] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[12][23] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[12][24] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[12][25] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[12][26] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[12][27] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[12][28] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[12][2] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[12][3] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[12][4] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[12][5] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[12][6] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[12][7] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[12][8] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[12][9] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[13][0] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[13][10] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[13][11] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[13][12] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[13][13] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[13][14] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[13][15] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[13][16] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[13][17] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[13][18] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[13][19] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[13][1] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[13][20] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[13][21] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[13][22] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[13][23] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[13][24] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[13][25] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[13][26] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[13][27] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[13][28] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[13][2] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[13][3] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[13][4] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[13][5] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[13][6] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[13][7] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[13][8] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[13][9] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[14][0] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[14][10] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[14][11] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[14][12] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[14][13] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[14][14] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[14][15] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[14][16] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[14][17] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[14][18] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[14][19] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[14][1] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[14][20] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[14][21] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[14][22] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[14][23] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[14][24] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[14][25] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[14][26] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[14][27] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[14][28] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[14][2] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[14][3] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[14][4] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[14][5] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[14][6] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[14][7] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[14][8] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[14][9] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[15][0] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[15][10] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[15][11] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[15][12] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[15][13] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[15][14] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[15][15] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[15][16] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[15][17] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[15][18] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[15][19] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[15][1] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[15][20] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[15][21] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[15][22] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[15][23] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[15][24] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[15][25] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[15][26] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[15][27] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[15][28] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[15][2] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[15][3] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[15][4] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[15][5] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[15][6] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[15][7] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[15][8] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[15][9] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[16][0] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[16][10] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[16][11] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[16][12] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[16][13] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[16][14] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[16][15] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[16][16] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[16][17] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[16][18] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[16][19] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[16][1] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[16][20] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[16][21] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[16][22] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[16][23] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[16][24] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[16][25] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[16][26] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[16][27] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[16][28] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[16][2] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[16][3] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[16][4] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[16][5] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[16][6] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[16][7] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[16][8] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[16][9] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[17][0] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[17][10] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[17][11] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[17][12] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[17][13] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[17][14] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[17][15] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[17][16] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[17][17] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[17][18] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[17][19] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[17][1] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[17][20] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[17][21] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[17][22] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[17][23] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[17][24] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[17][25] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[17][26] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[17][27] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[17][28] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[17][2] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[17][3] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[17][4] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[17][5] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[17][6] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[17][7] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[17][8] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[17][9] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[18][0] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[18][10] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[18][11] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[18][12] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[18][13] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[18][14] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[18][15] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[18][16] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[18][17] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[18][18] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[18][19] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[18][1] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[18][20] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[18][21] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[18][22] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[18][23] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[18][24] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[18][25] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[18][26] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[18][27] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[18][28] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[18][2] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[18][3] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[18][4] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[18][5] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[18][6] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[18][7] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[18][8] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[18][9] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[19][0] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[19][10] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[19][11] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[19][12] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[19][13] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[19][14] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[19][15] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[19][16] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[19][17] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[19][18] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[19][19] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[19][1] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[19][20] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[19][21] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[19][22] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[19][23] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[19][24] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[19][25] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[19][26] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[19][27] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[19][28] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[19][2] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[19][3] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[19][4] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[19][5] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[19][6] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[19][7] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[19][8] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[19][9] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[1][0] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[1][10] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[1][11] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[1][12] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[1][13] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[1][14] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[1][15] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[1][16] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[1][17] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[1][18] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[1][19] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[1][1] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[1][20] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[1][21] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[1][22] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[1][23] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[1][24] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[1][25] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[1][26] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[1][27] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[1][28] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[1][2] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[1][3] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[1][4] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[1][5] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[1][6] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[1][7] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[1][8] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[1][9] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[20][0] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[20][10] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[20][11] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[20][12] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[20][13] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[20][14] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[20][15] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[20][16] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[20][17] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[20][18] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[20][19] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[20][1] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[20][20] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[20][21] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[20][22] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[20][23] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[20][24] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[20][25] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[20][26] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[20][27] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[20][28] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[20][2] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[20][3] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[20][4] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[20][5] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[20][6] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[20][7] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[20][8] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[20][9] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[21][0] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[21][10] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[21][11] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[21][12] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[21][13] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[21][14] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[21][15] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[21][16] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[21][17] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[21][18] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[21][19] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[21][1] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[21][20] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[21][21] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[21][22] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[21][23] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[21][24] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[21][25] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[21][26] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[21][27] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[21][28] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[21][2] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[21][3] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[21][4] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[21][5] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[21][6] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[21][7] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[21][8] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[21][9] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[22][0] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[22][10] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[22][11] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[22][12] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[22][13] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[22][14] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[22][15] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[22][16] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[22][17] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[22][18] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[22][19] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[22][1] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[22][20] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[22][21] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[22][22] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[22][23] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[22][24] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[22][25] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[22][26] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[22][27] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[22][28] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[22][2] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[22][3] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[22][4] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[22][5] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[22][6] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[22][7] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[22][8] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[22][9] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[23][0] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[23][10] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[23][11] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[23][12] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[23][13] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[23][14] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[23][15] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[23][16] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[23][17] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[23][18] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[23][19] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[23][1] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[23][20] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[23][21] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[23][22] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[23][23] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[23][24] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[23][25] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[23][26] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[23][27] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[23][28] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[23][2] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[23][3] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[23][4] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[23][5] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[23][6] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[23][7] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[23][8] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[23][9] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[24][0] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[24][10] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[24][11] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[24][12] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[24][13] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[24][14] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[24][15] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[24][16] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[24][17] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[24][18] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[24][19] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[24][1] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[24][20] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[24][21] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[24][22] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[24][23] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[24][24] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[24][25] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[24][26] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[24][27] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[24][28] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[24][2] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[24][3] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[24][4] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[24][5] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[24][6] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[24][7] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[24][8] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[24][9] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[25][0] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[25][10] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[25][11] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[25][12] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[25][13] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[25][14] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[25][15] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[25][16] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[25][17] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[25][18] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[25][19] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[25][1] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[25][20] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[25][21] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[25][22] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[25][23] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[25][24] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[25][25] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[25][26] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[25][27] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[25][28] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[25][2] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[25][3] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[25][4] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[25][5] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[25][6] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[25][7] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[25][8] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[25][9] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[26][0] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[26][10] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[26][11] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[26][12] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[26][13] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[26][14] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[26][15] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[26][16] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[26][17] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[26][18] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[26][19] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[26][1] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[26][20] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[26][21] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[26][22] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[26][23] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[26][24] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[26][25] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[26][26] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[26][27] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[26][28] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[26][2] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[26][3] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[26][4] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[26][5] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[26][6] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[26][7] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[26][8] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[26][9] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[27][0] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[27][10] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[27][11] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[27][12] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[27][13] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[27][14] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[27][15] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[27][16] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[27][17] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[27][18] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[27][19] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[27][1] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[27][20] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[27][21] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[27][22] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[27][23] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[27][24] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[27][25] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[27][26] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[27][27] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[27][28] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[27][2] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[27][3] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[27][4] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[27][5] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[27][6] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[27][7] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[27][8] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[27][9] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[28][0] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[28][10] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[28][11] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[28][12] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[28][13] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[28][14] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[28][15] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[28][16] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[28][17] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[28][18] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[28][19] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[28][1] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[28][20] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[28][21] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[28][22] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[28][23] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[28][24] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[28][25] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[28][26] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[28][27] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[28][28] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[28][2] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[28][3] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[28][4] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[28][5] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[28][6] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[28][7] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[28][8] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[28][9] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[29][0] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[29][10] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[29][11] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[29][12] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[29][13] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[29][14] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[29][15] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[29][16] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[29][17] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[29][18] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[29][19] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[29][1] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[29][20] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[29][21] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[29][22] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[29][23] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[29][24] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[29][25] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[29][26] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[29][27] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[29][28] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[29][2] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[29][3] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[29][4] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[29][5] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[29][6] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[29][7] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[29][8] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[29][9] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[2][0] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[2][10] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[2][11] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[2][12] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[2][13] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[2][14] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[2][15] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[2][16] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[2][17] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[2][18] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[2][19] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[2][1] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[2][20] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[2][21] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[2][22] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[2][23] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[2][24] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[2][25] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[2][26] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[2][27] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[2][28] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[2][2] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[2][3] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[2][4] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[2][5] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[2][6] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[2][7] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[2][8] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[2][9] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[30][0] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[30][10] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[30][11] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[30][12] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[30][13] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[30][14] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[30][15] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[30][16] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[30][17] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[30][18] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[30][19] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[30][1] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[30][20] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[30][21] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[30][22] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[30][23] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[30][24] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[30][25] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[30][26] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[30][27] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[30][28] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[30][2] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[30][3] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[30][4] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[30][5] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[30][6] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[30][7] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[30][8] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[30][9] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[31][0] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[31][10] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[31][11] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[31][12] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[31][13] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[31][14] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[31][15] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[31][16] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[31][17] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[31][18] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[31][19] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[31][1] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[31][20] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[31][21] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[31][22] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[31][23] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[31][24] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[31][25] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[31][26] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[31][27] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[31][28] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[31][2] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[31][3] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[31][4] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[31][5] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[31][6] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[31][7] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[31][8] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[31][9] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[3][0] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[3][10] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[3][11] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[3][12] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[3][13] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[3][14] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[3][15] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[3][16] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[3][17] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[3][18] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[3][19] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[3][1] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[3][20] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[3][21] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[3][22] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[3][23] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[3][24] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[3][25] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[3][26] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[3][27] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[3][28] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[3][2] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[3][3] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[3][4] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[3][5] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[3][6] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[3][7] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[3][8] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[3][9] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[4][0] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[4][10] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[4][11] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[4][12] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[4][13] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[4][14] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[4][15] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[4][16] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[4][17] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[4][18] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[4][19] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[4][1] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[4][20] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[4][21] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[4][22] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[4][23] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[4][24] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[4][25] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[4][26] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[4][27] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[4][28] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[4][2] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[4][3] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[4][4] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[4][5] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[4][6] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[4][7] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[4][8] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[4][9] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[5][0] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[5][10] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[5][11] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[5][12] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[5][13] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[5][14] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[5][15] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[5][16] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[5][17] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[5][18] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[5][19] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[5][1] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[5][20] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[5][21] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[5][22] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[5][23] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[5][24] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[5][25] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[5][26] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[5][27] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[5][28] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[5][2] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[5][3] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[5][4] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[5][5] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[5][6] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[5][7] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[5][8] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[5][9] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[6][0] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[6][10] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[6][11] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[6][12] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[6][13] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[6][14] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[6][15] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[6][16] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[6][17] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[6][18] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[6][19] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[6][1] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[6][20] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[6][21] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[6][22] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[6][23] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[6][24] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[6][25] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[6][26] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[6][27] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[6][28] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[6][2] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[6][3] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[6][4] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[6][5] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[6][6] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[6][7] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[6][8] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[6][9] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[7][0] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[7][10] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[7][11] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[7][12] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[7][13] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[7][14] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[7][15] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[7][16] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[7][17] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[7][18] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[7][19] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[7][1] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[7][20] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[7][21] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[7][22] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[7][23] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[7][24] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[7][25] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[7][26] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[7][27] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[7][28] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[7][2] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[7][3] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[7][4] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[7][5] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[7][6] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[7][7] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[7][8] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[7][9] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[8][0] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[8][10] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[8][11] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[8][12] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[8][13] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[8][14] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[8][15] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[8][16] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[8][17] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[8][18] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[8][19] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[8][1] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[8][20] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[8][21] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[8][22] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[8][23] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[8][24] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[8][25] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[8][26] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[8][27] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[8][28] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[8][2] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[8][3] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[8][4] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[8][5] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[8][6] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[8][7] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[8][8] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[8][9] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[9][0] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[9][10] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[9][11] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[9][12] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[9][13] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[9][14] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[9][15] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[9][16] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[9][17] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[9][18] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[9][19] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[9][1] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[9][20] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[9][21] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[9][22] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[9][23] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[9][24] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[9][25] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[9][26] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[9][27] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[9][28] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[9][2] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[9][3] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[9][4] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[9][5] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[9][6] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[9][7] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[9][8] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[9][9] ;
 wire \soc.spi_video_ram_1.write_fifo.read_pointer[0] ;
 wire \soc.spi_video_ram_1.write_fifo.read_pointer[1] ;
 wire \soc.spi_video_ram_1.write_fifo.read_pointer[2] ;
 wire \soc.spi_video_ram_1.write_fifo.read_pointer[3] ;
 wire \soc.spi_video_ram_1.write_fifo.read_pointer[4] ;
 wire \soc.spi_video_ram_1.write_fifo.write_pointer[0] ;
 wire \soc.spi_video_ram_1.write_fifo.write_pointer[1] ;
 wire \soc.spi_video_ram_1.write_fifo.write_pointer[2] ;
 wire \soc.spi_video_ram_1.write_fifo.write_pointer[3] ;
 wire \soc.spi_video_ram_1.write_fifo.write_pointer[4] ;
 wire \soc.synch_hack_writeM ;
 wire \soc.video_generator_1.h_count[1] ;
 wire \soc.video_generator_1.h_count[2] ;
 wire \soc.video_generator_1.h_count[3] ;
 wire \soc.video_generator_1.h_count[4] ;
 wire \soc.video_generator_1.h_count[5] ;
 wire \soc.video_generator_1.h_count[6] ;
 wire \soc.video_generator_1.h_count[7] ;
 wire \soc.video_generator_1.h_count[8] ;
 wire \soc.video_generator_1.h_count[9] ;
 wire \soc.video_generator_1.v_count[0] ;
 wire \soc.video_generator_1.v_count[1] ;
 wire \soc.video_generator_1.v_count[2] ;
 wire \soc.video_generator_1.v_count[3] ;
 wire \soc.video_generator_1.v_count[4] ;
 wire \soc.video_generator_1.v_count[5] ;
 wire \soc.video_generator_1.v_count[6] ;
 wire \soc.video_generator_1.v_count[7] ;
 wire \soc.video_generator_1.v_count[8] ;
 wire \soc.video_generator_1.v_count[9] ;
 wire net192;
 wire net193;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net194;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net195;
 wire net223;
 wire net224;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire clknet_leaf_1_wb_clk_i;
 wire clknet_leaf_2_wb_clk_i;
 wire clknet_leaf_3_wb_clk_i;
 wire clknet_leaf_4_wb_clk_i;
 wire clknet_leaf_5_wb_clk_i;
 wire clknet_leaf_6_wb_clk_i;
 wire clknet_leaf_7_wb_clk_i;
 wire clknet_leaf_8_wb_clk_i;
 wire clknet_leaf_9_wb_clk_i;
 wire clknet_leaf_10_wb_clk_i;
 wire clknet_leaf_11_wb_clk_i;
 wire clknet_leaf_12_wb_clk_i;
 wire clknet_leaf_13_wb_clk_i;
 wire clknet_leaf_14_wb_clk_i;
 wire clknet_leaf_15_wb_clk_i;
 wire clknet_leaf_16_wb_clk_i;
 wire clknet_leaf_17_wb_clk_i;
 wire clknet_leaf_18_wb_clk_i;
 wire clknet_leaf_19_wb_clk_i;
 wire clknet_leaf_20_wb_clk_i;
 wire clknet_leaf_21_wb_clk_i;
 wire clknet_leaf_22_wb_clk_i;
 wire clknet_leaf_23_wb_clk_i;
 wire clknet_leaf_24_wb_clk_i;
 wire clknet_leaf_25_wb_clk_i;
 wire clknet_leaf_26_wb_clk_i;
 wire clknet_leaf_27_wb_clk_i;
 wire clknet_leaf_28_wb_clk_i;
 wire clknet_leaf_29_wb_clk_i;
 wire clknet_leaf_30_wb_clk_i;
 wire clknet_leaf_31_wb_clk_i;
 wire clknet_leaf_32_wb_clk_i;
 wire clknet_leaf_33_wb_clk_i;
 wire clknet_leaf_34_wb_clk_i;
 wire clknet_leaf_35_wb_clk_i;
 wire clknet_leaf_36_wb_clk_i;
 wire clknet_leaf_37_wb_clk_i;
 wire clknet_leaf_38_wb_clk_i;
 wire clknet_leaf_39_wb_clk_i;
 wire clknet_leaf_40_wb_clk_i;
 wire clknet_leaf_41_wb_clk_i;
 wire clknet_leaf_42_wb_clk_i;
 wire clknet_leaf_43_wb_clk_i;
 wire clknet_leaf_44_wb_clk_i;
 wire clknet_leaf_45_wb_clk_i;
 wire clknet_leaf_46_wb_clk_i;
 wire clknet_leaf_47_wb_clk_i;
 wire clknet_leaf_48_wb_clk_i;
 wire clknet_leaf_49_wb_clk_i;
 wire clknet_leaf_50_wb_clk_i;
 wire clknet_leaf_51_wb_clk_i;
 wire clknet_leaf_52_wb_clk_i;
 wire clknet_leaf_53_wb_clk_i;
 wire clknet_leaf_54_wb_clk_i;
 wire clknet_leaf_55_wb_clk_i;
 wire clknet_leaf_56_wb_clk_i;
 wire clknet_leaf_58_wb_clk_i;
 wire clknet_leaf_59_wb_clk_i;
 wire clknet_leaf_60_wb_clk_i;
 wire clknet_leaf_61_wb_clk_i;
 wire clknet_leaf_62_wb_clk_i;
 wire clknet_leaf_63_wb_clk_i;
 wire clknet_leaf_64_wb_clk_i;
 wire clknet_leaf_65_wb_clk_i;
 wire clknet_leaf_66_wb_clk_i;
 wire clknet_leaf_67_wb_clk_i;
 wire clknet_leaf_68_wb_clk_i;
 wire clknet_leaf_69_wb_clk_i;
 wire clknet_leaf_70_wb_clk_i;
 wire clknet_leaf_71_wb_clk_i;
 wire clknet_leaf_72_wb_clk_i;
 wire clknet_leaf_73_wb_clk_i;
 wire clknet_leaf_74_wb_clk_i;
 wire clknet_leaf_75_wb_clk_i;
 wire clknet_leaf_76_wb_clk_i;
 wire clknet_leaf_77_wb_clk_i;
 wire clknet_leaf_78_wb_clk_i;
 wire clknet_leaf_79_wb_clk_i;
 wire clknet_leaf_80_wb_clk_i;
 wire clknet_leaf_81_wb_clk_i;
 wire clknet_leaf_82_wb_clk_i;
 wire clknet_leaf_83_wb_clk_i;
 wire clknet_leaf_85_wb_clk_i;
 wire clknet_leaf_86_wb_clk_i;
 wire clknet_leaf_87_wb_clk_i;
 wire clknet_leaf_89_wb_clk_i;
 wire clknet_leaf_92_wb_clk_i;
 wire clknet_leaf_93_wb_clk_i;
 wire clknet_leaf_95_wb_clk_i;
 wire clknet_leaf_96_wb_clk_i;
 wire clknet_leaf_97_wb_clk_i;
 wire clknet_leaf_98_wb_clk_i;
 wire clknet_leaf_99_wb_clk_i;
 wire clknet_leaf_100_wb_clk_i;
 wire clknet_leaf_101_wb_clk_i;
 wire clknet_leaf_102_wb_clk_i;
 wire clknet_leaf_104_wb_clk_i;
 wire clknet_leaf_105_wb_clk_i;
 wire clknet_leaf_106_wb_clk_i;
 wire clknet_leaf_107_wb_clk_i;
 wire clknet_leaf_108_wb_clk_i;
 wire clknet_leaf_109_wb_clk_i;
 wire clknet_leaf_110_wb_clk_i;
 wire clknet_leaf_111_wb_clk_i;
 wire clknet_leaf_112_wb_clk_i;
 wire clknet_leaf_113_wb_clk_i;
 wire clknet_leaf_114_wb_clk_i;
 wire clknet_leaf_115_wb_clk_i;
 wire clknet_leaf_117_wb_clk_i;
 wire clknet_leaf_118_wb_clk_i;
 wire clknet_leaf_119_wb_clk_i;
 wire clknet_leaf_121_wb_clk_i;
 wire clknet_leaf_122_wb_clk_i;
 wire clknet_leaf_123_wb_clk_i;
 wire clknet_leaf_124_wb_clk_i;
 wire clknet_leaf_125_wb_clk_i;
 wire clknet_leaf_126_wb_clk_i;
 wire clknet_leaf_127_wb_clk_i;
 wire clknet_leaf_128_wb_clk_i;
 wire clknet_leaf_129_wb_clk_i;
 wire clknet_leaf_130_wb_clk_i;
 wire clknet_leaf_132_wb_clk_i;
 wire clknet_leaf_134_wb_clk_i;
 wire clknet_leaf_135_wb_clk_i;
 wire clknet_leaf_136_wb_clk_i;
 wire clknet_leaf_137_wb_clk_i;
 wire clknet_leaf_138_wb_clk_i;
 wire clknet_leaf_139_wb_clk_i;
 wire clknet_leaf_140_wb_clk_i;
 wire clknet_leaf_141_wb_clk_i;
 wire clknet_leaf_142_wb_clk_i;
 wire clknet_leaf_143_wb_clk_i;
 wire clknet_leaf_144_wb_clk_i;
 wire clknet_leaf_145_wb_clk_i;
 wire clknet_leaf_146_wb_clk_i;
 wire clknet_leaf_147_wb_clk_i;
 wire clknet_leaf_148_wb_clk_i;
 wire clknet_leaf_149_wb_clk_i;
 wire clknet_leaf_150_wb_clk_i;
 wire clknet_leaf_151_wb_clk_i;
 wire clknet_leaf_152_wb_clk_i;
 wire clknet_leaf_153_wb_clk_i;
 wire clknet_leaf_154_wb_clk_i;
 wire clknet_leaf_155_wb_clk_i;
 wire clknet_leaf_156_wb_clk_i;
 wire clknet_leaf_157_wb_clk_i;
 wire clknet_leaf_158_wb_clk_i;
 wire clknet_leaf_159_wb_clk_i;
 wire clknet_leaf_160_wb_clk_i;
 wire clknet_leaf_161_wb_clk_i;
 wire clknet_leaf_162_wb_clk_i;
 wire clknet_leaf_163_wb_clk_i;
 wire clknet_leaf_164_wb_clk_i;
 wire clknet_leaf_165_wb_clk_i;
 wire clknet_leaf_166_wb_clk_i;
 wire clknet_leaf_167_wb_clk_i;
 wire clknet_leaf_168_wb_clk_i;
 wire clknet_leaf_169_wb_clk_i;
 wire clknet_leaf_170_wb_clk_i;
 wire clknet_leaf_173_wb_clk_i;
 wire clknet_leaf_175_wb_clk_i;
 wire clknet_leaf_176_wb_clk_i;
 wire clknet_leaf_177_wb_clk_i;
 wire clknet_leaf_178_wb_clk_i;
 wire clknet_leaf_179_wb_clk_i;
 wire clknet_leaf_180_wb_clk_i;
 wire clknet_leaf_183_wb_clk_i;
 wire clknet_leaf_184_wb_clk_i;
 wire clknet_leaf_185_wb_clk_i;
 wire clknet_leaf_186_wb_clk_i;
 wire clknet_leaf_187_wb_clk_i;
 wire clknet_leaf_188_wb_clk_i;
 wire clknet_leaf_189_wb_clk_i;
 wire clknet_leaf_190_wb_clk_i;
 wire clknet_leaf_191_wb_clk_i;
 wire clknet_leaf_192_wb_clk_i;
 wire clknet_leaf_193_wb_clk_i;
 wire clknet_leaf_194_wb_clk_i;
 wire clknet_leaf_195_wb_clk_i;
 wire clknet_leaf_196_wb_clk_i;
 wire clknet_leaf_197_wb_clk_i;
 wire clknet_leaf_198_wb_clk_i;
 wire clknet_leaf_199_wb_clk_i;
 wire clknet_leaf_200_wb_clk_i;
 wire clknet_leaf_201_wb_clk_i;
 wire clknet_leaf_202_wb_clk_i;
 wire clknet_leaf_203_wb_clk_i;
 wire clknet_leaf_205_wb_clk_i;
 wire clknet_leaf_207_wb_clk_i;
 wire clknet_leaf_208_wb_clk_i;
 wire clknet_leaf_210_wb_clk_i;
 wire clknet_leaf_211_wb_clk_i;
 wire clknet_leaf_212_wb_clk_i;
 wire clknet_leaf_213_wb_clk_i;
 wire clknet_leaf_214_wb_clk_i;
 wire clknet_leaf_215_wb_clk_i;
 wire clknet_leaf_216_wb_clk_i;
 wire clknet_leaf_217_wb_clk_i;
 wire clknet_leaf_218_wb_clk_i;
 wire clknet_leaf_219_wb_clk_i;
 wire clknet_leaf_220_wb_clk_i;
 wire clknet_leaf_221_wb_clk_i;
 wire clknet_leaf_222_wb_clk_i;
 wire clknet_leaf_224_wb_clk_i;
 wire clknet_leaf_226_wb_clk_i;
 wire clknet_leaf_227_wb_clk_i;
 wire clknet_leaf_228_wb_clk_i;
 wire clknet_leaf_229_wb_clk_i;
 wire clknet_leaf_230_wb_clk_i;
 wire clknet_leaf_231_wb_clk_i;
 wire clknet_leaf_232_wb_clk_i;
 wire clknet_leaf_233_wb_clk_i;
 wire clknet_leaf_234_wb_clk_i;
 wire clknet_leaf_235_wb_clk_i;
 wire clknet_leaf_236_wb_clk_i;
 wire clknet_leaf_237_wb_clk_i;
 wire clknet_leaf_238_wb_clk_i;
 wire clknet_leaf_239_wb_clk_i;
 wire clknet_leaf_240_wb_clk_i;
 wire clknet_leaf_241_wb_clk_i;
 wire clknet_leaf_242_wb_clk_i;
 wire clknet_leaf_243_wb_clk_i;
 wire clknet_leaf_244_wb_clk_i;
 wire clknet_leaf_245_wb_clk_i;
 wire clknet_leaf_246_wb_clk_i;
 wire clknet_leaf_247_wb_clk_i;
 wire clknet_leaf_248_wb_clk_i;
 wire clknet_leaf_249_wb_clk_i;
 wire clknet_leaf_250_wb_clk_i;
 wire clknet_leaf_251_wb_clk_i;
 wire clknet_leaf_252_wb_clk_i;
 wire clknet_leaf_253_wb_clk_i;
 wire clknet_leaf_254_wb_clk_i;
 wire clknet_leaf_255_wb_clk_i;
 wire clknet_leaf_256_wb_clk_i;
 wire clknet_leaf_257_wb_clk_i;
 wire clknet_leaf_258_wb_clk_i;
 wire clknet_leaf_259_wb_clk_i;
 wire clknet_leaf_260_wb_clk_i;
 wire clknet_leaf_261_wb_clk_i;
 wire clknet_leaf_262_wb_clk_i;
 wire clknet_leaf_263_wb_clk_i;
 wire clknet_leaf_264_wb_clk_i;
 wire clknet_leaf_265_wb_clk_i;
 wire clknet_leaf_266_wb_clk_i;
 wire clknet_leaf_267_wb_clk_i;
 wire clknet_leaf_268_wb_clk_i;
 wire clknet_leaf_269_wb_clk_i;
 wire clknet_leaf_270_wb_clk_i;
 wire clknet_leaf_271_wb_clk_i;
 wire clknet_leaf_272_wb_clk_i;
 wire clknet_leaf_273_wb_clk_i;
 wire clknet_leaf_274_wb_clk_i;
 wire clknet_leaf_276_wb_clk_i;
 wire clknet_leaf_277_wb_clk_i;
 wire clknet_leaf_278_wb_clk_i;
 wire clknet_leaf_279_wb_clk_i;
 wire clknet_leaf_280_wb_clk_i;
 wire clknet_leaf_281_wb_clk_i;
 wire clknet_leaf_282_wb_clk_i;
 wire clknet_leaf_283_wb_clk_i;
 wire clknet_leaf_284_wb_clk_i;
 wire clknet_leaf_285_wb_clk_i;
 wire clknet_leaf_286_wb_clk_i;
 wire clknet_leaf_287_wb_clk_i;
 wire clknet_leaf_288_wb_clk_i;
 wire clknet_leaf_289_wb_clk_i;
 wire clknet_leaf_290_wb_clk_i;
 wire clknet_leaf_291_wb_clk_i;
 wire clknet_leaf_292_wb_clk_i;
 wire clknet_leaf_293_wb_clk_i;
 wire clknet_leaf_294_wb_clk_i;
 wire clknet_leaf_295_wb_clk_i;
 wire clknet_leaf_296_wb_clk_i;
 wire clknet_leaf_297_wb_clk_i;
 wire clknet_leaf_298_wb_clk_i;
 wire clknet_leaf_299_wb_clk_i;
 wire clknet_leaf_300_wb_clk_i;
 wire clknet_leaf_301_wb_clk_i;
 wire clknet_leaf_302_wb_clk_i;
 wire clknet_leaf_303_wb_clk_i;
 wire clknet_leaf_304_wb_clk_i;
 wire clknet_leaf_305_wb_clk_i;
 wire clknet_leaf_306_wb_clk_i;
 wire clknet_leaf_307_wb_clk_i;
 wire clknet_leaf_308_wb_clk_i;
 wire clknet_leaf_309_wb_clk_i;
 wire clknet_leaf_310_wb_clk_i;
 wire clknet_leaf_311_wb_clk_i;
 wire clknet_leaf_312_wb_clk_i;
 wire clknet_leaf_313_wb_clk_i;
 wire clknet_leaf_314_wb_clk_i;
 wire clknet_leaf_315_wb_clk_i;
 wire clknet_leaf_316_wb_clk_i;
 wire clknet_leaf_317_wb_clk_i;
 wire clknet_leaf_318_wb_clk_i;
 wire clknet_leaf_319_wb_clk_i;
 wire clknet_leaf_320_wb_clk_i;
 wire clknet_leaf_321_wb_clk_i;
 wire clknet_0_wb_clk_i;
 wire clknet_2_0_0_wb_clk_i;
 wire clknet_2_1_0_wb_clk_i;
 wire clknet_2_2_0_wb_clk_i;
 wire clknet_2_3_0_wb_clk_i;
 wire clknet_3_0_0_wb_clk_i;
 wire clknet_3_1_0_wb_clk_i;
 wire clknet_3_2_0_wb_clk_i;
 wire clknet_3_3_0_wb_clk_i;
 wire clknet_3_4_0_wb_clk_i;
 wire clknet_3_5_0_wb_clk_i;
 wire clknet_3_6_0_wb_clk_i;
 wire clknet_3_7_0_wb_clk_i;
 wire clknet_4_0_0_wb_clk_i;
 wire clknet_4_1_0_wb_clk_i;
 wire clknet_4_2_0_wb_clk_i;
 wire clknet_4_3_0_wb_clk_i;
 wire clknet_4_4_0_wb_clk_i;
 wire clknet_4_5_0_wb_clk_i;
 wire clknet_4_6_0_wb_clk_i;
 wire clknet_4_7_0_wb_clk_i;
 wire clknet_4_8_0_wb_clk_i;
 wire clknet_4_9_0_wb_clk_i;
 wire clknet_4_10_0_wb_clk_i;
 wire clknet_4_11_0_wb_clk_i;
 wire clknet_4_12_0_wb_clk_i;
 wire clknet_4_13_0_wb_clk_i;
 wire clknet_4_14_0_wb_clk_i;
 wire clknet_4_15_0_wb_clk_i;
 wire clknet_5_0_0_wb_clk_i;
 wire clknet_5_1_0_wb_clk_i;
 wire clknet_5_2_0_wb_clk_i;
 wire clknet_5_3_0_wb_clk_i;
 wire clknet_5_4_0_wb_clk_i;
 wire clknet_5_5_0_wb_clk_i;
 wire clknet_5_6_0_wb_clk_i;
 wire clknet_5_7_0_wb_clk_i;
 wire clknet_5_8_0_wb_clk_i;
 wire clknet_5_9_0_wb_clk_i;
 wire clknet_5_10_0_wb_clk_i;
 wire clknet_5_11_0_wb_clk_i;
 wire clknet_5_12_0_wb_clk_i;
 wire clknet_5_13_0_wb_clk_i;
 wire clknet_5_14_0_wb_clk_i;
 wire clknet_5_15_0_wb_clk_i;
 wire clknet_5_16_0_wb_clk_i;
 wire clknet_5_17_0_wb_clk_i;
 wire clknet_5_18_0_wb_clk_i;
 wire clknet_5_19_0_wb_clk_i;
 wire clknet_5_20_0_wb_clk_i;
 wire clknet_5_21_0_wb_clk_i;
 wire clknet_5_22_0_wb_clk_i;
 wire clknet_5_23_0_wb_clk_i;
 wire clknet_5_24_0_wb_clk_i;
 wire clknet_5_25_0_wb_clk_i;
 wire clknet_5_26_0_wb_clk_i;
 wire clknet_5_27_0_wb_clk_i;
 wire clknet_5_28_0_wb_clk_i;
 wire clknet_5_29_0_wb_clk_i;
 wire clknet_5_30_0_wb_clk_i;
 wire clknet_5_31_0_wb_clk_i;
 wire clknet_opt_1_0_wb_clk_i;
 wire clknet_opt_2_0_wb_clk_i;
 wire clknet_opt_3_0_wb_clk_i;
 wire clknet_opt_4_0_wb_clk_i;
 wire clknet_opt_5_0_wb_clk_i;

 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 _05462_ (.I(net18),
    .Z(_01378_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_4 _05463_ (.I(_01378_),
    .ZN(_01379_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 _05464_ (.I(_01379_),
    .Z(_01380_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05465_ (.I(_01380_),
    .Z(_01381_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _05466_ (.A1(\soc.spi_video_ram_1.state_counter[9] ),
    .A2(\soc.spi_video_ram_1.state_counter[8] ),
    .A3(\soc.spi_video_ram_1.state_counter[10] ),
    .ZN(_01382_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _05467_ (.A1(\soc.spi_video_ram_1.state_counter[5] ),
    .A2(\soc.spi_video_ram_1.state_counter[4] ),
    .A3(\soc.spi_video_ram_1.state_counter[7] ),
    .A4(\soc.spi_video_ram_1.state_counter[6] ),
    .ZN(_01383_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _05468_ (.A1(\soc.spi_video_ram_1.state_counter[1] ),
    .A2(\soc.spi_video_ram_1.state_counter[0] ),
    .A3(\soc.spi_video_ram_1.state_counter[3] ),
    .A4(\soc.spi_video_ram_1.state_counter[2] ),
    .ZN(_01384_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _05469_ (.A1(_01382_),
    .A2(_01383_),
    .A3(_01384_),
    .ZN(_01385_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _05470_ (.I(\soc.spi_video_ram_1.state_sram_clk_counter[1] ),
    .ZN(_01386_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _05471_ (.I(\soc.spi_video_ram_1.state_sram_clk_counter[8] ),
    .Z(_01387_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _05472_ (.A1(\soc.spi_video_ram_1.state_sram_clk_counter[7] ),
    .A2(\soc.spi_video_ram_1.state_sram_clk_counter[6] ),
    .A3(\soc.spi_video_ram_1.state_sram_clk_counter[5] ),
    .A4(\soc.spi_video_ram_1.state_sram_clk_counter[4] ),
    .ZN(_01388_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05473_ (.A1(\soc.spi_video_ram_1.state_sram_clk_counter[3] ),
    .A2(\soc.spi_video_ram_1.state_sram_clk_counter[2] ),
    .ZN(_01389_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05474_ (.A1(_01388_),
    .A2(_01389_),
    .ZN(_01390_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _05475_ (.A1(_01387_),
    .A2(\soc.spi_video_ram_1.state_sram_clk_counter[0] ),
    .A3(_01390_),
    .Z(_01391_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _05476_ (.A1(_01386_),
    .A2(_01391_),
    .ZN(_01392_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05477_ (.A1(_01385_),
    .A2(_01392_),
    .ZN(_01393_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05478_ (.A1(\soc.spi_video_ram_1.current_state[0] ),
    .A2(_01393_),
    .ZN(_01394_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05479_ (.A1(_01381_),
    .A2(_01394_),
    .ZN(_00005_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05480_ (.I(_01378_),
    .Z(_01395_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05481_ (.I(_01395_),
    .Z(_01396_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05482_ (.I(_01393_),
    .ZN(_01397_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _05483_ (.A1(\soc.spi_video_ram_1.write_fifo.read_pointer[2] ),
    .A2(\soc.spi_video_ram_1.write_fifo.write_pointer[2] ),
    .Z(_01398_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05484_ (.I(_01398_),
    .ZN(_01399_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _05485_ (.I(\soc.spi_video_ram_1.write_fifo.write_pointer[1] ),
    .ZN(_01400_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _05486_ (.A1(\soc.spi_video_ram_1.write_fifo.read_pointer[1] ),
    .A2(_01400_),
    .Z(_01401_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05487_ (.A1(_01399_),
    .A2(_01401_),
    .ZN(_01402_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 _05488_ (.I(\soc.spi_video_ram_1.write_fifo.write_pointer[3] ),
    .Z(_01403_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _05489_ (.A1(\soc.spi_video_ram_1.write_fifo.read_pointer[3] ),
    .A2(_01403_),
    .Z(_01404_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 _05490_ (.I(\soc.spi_video_ram_1.write_fifo.write_pointer[0] ),
    .Z(_01405_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _05491_ (.A1(\soc.spi_video_ram_1.write_fifo.read_pointer[0] ),
    .A2(_01405_),
    .Z(_01406_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _05492_ (.A1(\soc.spi_video_ram_1.write_fifo.read_pointer[4] ),
    .A2(\soc.spi_video_ram_1.write_fifo.write_pointer[4] ),
    .Z(_01407_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _05493_ (.A1(_01402_),
    .A2(_01404_),
    .A3(_01406_),
    .A4(_01407_),
    .ZN(_01408_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05494_ (.I(\soc.spi_video_ram_1.current_state[3] ),
    .ZN(_01409_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05495_ (.A1(\soc.spi_video_ram_1.current_state[1] ),
    .A2(\soc.spi_video_ram_1.current_state[4] ),
    .ZN(_01410_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _05496_ (.A1(_01409_),
    .A2(_01410_),
    .ZN(_01411_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _05497_ (.A1(\soc.spi_video_ram_1.current_state[0] ),
    .A2(_01408_),
    .A3(_01411_),
    .ZN(_01412_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05498_ (.A1(\soc.spi_video_ram_1.initialized ),
    .A2(\soc.spi_video_ram_1.current_state[2] ),
    .ZN(_01413_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _05499_ (.A1(\soc.spi_video_ram_1.start_read ),
    .A2(_01408_),
    .B(_01412_),
    .C(_01413_),
    .ZN(_01414_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05500_ (.I(\soc.spi_video_ram_1.state_sram_clk_counter[2] ),
    .ZN(_01415_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _05501_ (.A1(_01387_),
    .A2(\soc.spi_video_ram_1.state_sram_clk_counter[1] ),
    .A3(\soc.spi_video_ram_1.state_sram_clk_counter[0] ),
    .ZN(_01416_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _05502_ (.A1(\soc.spi_video_ram_1.state_sram_clk_counter[3] ),
    .A2(_01415_),
    .A3(_01388_),
    .A4(_01416_),
    .ZN(_01417_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _05503_ (.A1(_01409_),
    .A2(_01417_),
    .Z(_01418_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _05504_ (.I(\soc.spi_video_ram_1.current_state[4] ),
    .Z(_01419_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05505_ (.I(_01387_),
    .ZN(_01420_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _05506_ (.A1(\soc.spi_video_ram_1.state_sram_clk_counter[3] ),
    .A2(_01415_),
    .A3(\soc.spi_video_ram_1.state_sram_clk_counter[0] ),
    .Z(_01421_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _05507_ (.A1(_01420_),
    .A2(\soc.spi_video_ram_1.state_sram_clk_counter[7] ),
    .A3(\soc.spi_video_ram_1.state_sram_clk_counter[1] ),
    .A4(_01421_),
    .ZN(_01422_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _05508_ (.A1(\soc.spi_video_ram_1.state_sram_clk_counter[6] ),
    .A2(\soc.spi_video_ram_1.state_sram_clk_counter[5] ),
    .A3(\soc.spi_video_ram_1.state_sram_clk_counter[4] ),
    .A4(_01422_),
    .ZN(_01423_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _05509_ (.A1(\soc.spi_video_ram_1.state_sram_clk_counter[3] ),
    .A2(\soc.spi_video_ram_1.state_sram_clk_counter[2] ),
    .A3(_01388_),
    .A4(_01416_),
    .Z(_01424_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _05510_ (.A1(_01419_),
    .A2(_01423_),
    .B1(_01424_),
    .B2(\soc.spi_video_ram_1.current_state[1] ),
    .ZN(_01425_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05511_ (.A1(_01418_),
    .A2(_01425_),
    .ZN(_01426_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _05512_ (.A1(\soc.spi_video_ram_1.current_state[0] ),
    .A2(_01397_),
    .B(_01414_),
    .C(_01426_),
    .ZN(_01427_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05513_ (.A1(_01396_),
    .A2(_01427_),
    .ZN(_00007_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05514_ (.I(\soc.spi_video_ram_1.current_state[3] ),
    .Z(_01428_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05515_ (.A1(_01428_),
    .A2(_01417_),
    .ZN(_01429_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05516_ (.I(\soc.spi_video_ram_1.initialized ),
    .ZN(_01430_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05517_ (.A1(_01430_),
    .A2(\soc.spi_video_ram_1.current_state[2] ),
    .ZN(_01431_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05518_ (.A1(_01429_),
    .A2(_01431_),
    .B(_01396_),
    .ZN(_00008_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05519_ (.I(\soc.spi_video_ram_1.state_sram_clk_counter[7] ),
    .ZN(_01432_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _05520_ (.A1(_01432_),
    .A2(\soc.spi_video_ram_1.state_sram_clk_counter[6] ),
    .A3(\soc.spi_video_ram_1.state_sram_clk_counter[5] ),
    .A4(\soc.spi_video_ram_1.state_sram_clk_counter[4] ),
    .ZN(_01433_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _05521_ (.A1(_01420_),
    .A2(\soc.spi_video_ram_1.state_sram_clk_counter[1] ),
    .A3(_01421_),
    .A4(_01433_),
    .ZN(_01434_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05522_ (.A1(_01419_),
    .A2(_01434_),
    .ZN(_01435_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _05523_ (.A1(\soc.spi_video_ram_1.initialized ),
    .A2(\soc.spi_video_ram_1.start_read ),
    .A3(\soc.spi_video_ram_1.current_state[2] ),
    .A4(_01408_),
    .ZN(_01436_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05524_ (.A1(_01435_),
    .A2(_01436_),
    .B(_01396_),
    .ZN(_00009_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05525_ (.I(\soc.spi_video_ram_1.current_state[1] ),
    .ZN(_01437_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _05526_ (.A1(_01437_),
    .A2(_01424_),
    .Z(_01438_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _05527_ (.A1(\soc.spi_video_ram_1.current_state[2] ),
    .A2(_01412_),
    .Z(_01439_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05528_ (.I(_01439_),
    .Z(_00010_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05529_ (.A1(\soc.spi_video_ram_1.initialized ),
    .A2(_00010_),
    .ZN(_01440_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05530_ (.A1(_01438_),
    .A2(_01440_),
    .B(_01396_),
    .ZN(_00006_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _05531_ (.A1(\soc.spi_video_ram_1.write_fifo.write_pointer[1] ),
    .A2(_01405_),
    .ZN(_01441_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _05532_ (.A1(_01405_),
    .A2(_01401_),
    .B1(_01441_),
    .B2(_01398_),
    .ZN(_01442_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05533_ (.A1(_01405_),
    .A2(_01401_),
    .B(_01442_),
    .ZN(_01443_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _05534_ (.I(_01405_),
    .ZN(_01444_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _05535_ (.A1(_01400_),
    .A2(_01444_),
    .ZN(_01445_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05536_ (.A1(\soc.spi_video_ram_1.write_fifo.write_pointer[2] ),
    .A2(_01445_),
    .ZN(_01446_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _05537_ (.A1(_01404_),
    .A2(_01446_),
    .ZN(_01447_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05538_ (.A1(_01398_),
    .A2(_01441_),
    .B(_01447_),
    .ZN(_01448_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _05539_ (.A1(_01403_),
    .A2(\soc.spi_video_ram_1.write_fifo.write_pointer[2] ),
    .A3(_01445_),
    .ZN(_01449_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _05540_ (.A1(_01407_),
    .A2(_01449_),
    .Z(_01450_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _05541_ (.A1(_01406_),
    .A2(_01443_),
    .A3(_01448_),
    .A4(_01450_),
    .Z(_01451_));
 gf180mcu_fd_sc_mcu7t5v0__or4_2 _05542_ (.A1(\soc.rom_encoder_0.write_enable ),
    .A2(net18),
    .A3(net13),
    .A4(net37),
    .Z(_01452_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _05543_ (.A1(\soc.ram_encoder_0.initialized ),
    .A2(\soc.rom_encoder_0.initialized ),
    .A3(\soc.spi_video_ram_1.initialized ),
    .ZN(_01453_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _05544_ (.A1(\soc.hack_wait_clocks[1] ),
    .A2(\soc.hack_wait_clocks[0] ),
    .A3(_01452_),
    .A4(_01453_),
    .Z(_01454_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _05545_ (.A1(\soc.cpu.instruction[15] ),
    .A2(\soc.cpu.instruction[3] ),
    .ZN(_01455_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05546_ (.I(\soc.cpu.AReg.data[13] ),
    .ZN(_01456_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _05547_ (.A1(net87),
    .A2(\soc.hack_clk_strobe ),
    .A3(\soc.cpu.AReg.data[14] ),
    .A4(_01456_),
    .ZN(_01457_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _05548_ (.A1(_01451_),
    .A2(_01454_),
    .A3(_01455_),
    .A4(_01457_),
    .ZN(_01458_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 _05549_ (.I(_01458_),
    .Z(_01459_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05550_ (.I(_01459_),
    .Z(_00011_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _05551_ (.I(\soc.spi_video_ram_1.buffer_index[4] ),
    .ZN(_01460_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _05552_ (.I(\soc.spi_video_ram_1.buffer_index[0] ),
    .Z(_01461_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05553_ (.A1(_01461_),
    .A2(\soc.spi_video_ram_1.buffer_index[1] ),
    .ZN(_01462_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05554_ (.I(\soc.spi_video_ram_1.buffer_index[3] ),
    .Z(_01463_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _05555_ (.A1(\soc.spi_video_ram_1.buffer_index[2] ),
    .A2(_01463_),
    .ZN(_01464_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _05556_ (.A1(\soc.spi_video_ram_1.buffer_index[4] ),
    .A2(_01464_),
    .Z(_01465_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05557_ (.A1(_01462_),
    .A2(_01465_),
    .ZN(_01466_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05558_ (.I(_01461_),
    .Z(_01467_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 _05559_ (.I(_01467_),
    .Z(_01468_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05560_ (.I(\soc.spi_video_ram_1.buffer_index[1] ),
    .Z(_01469_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05561_ (.I(\soc.spi_video_ram_1.buffer_index[2] ),
    .Z(_01470_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _05562_ (.A1(_01469_),
    .A2(_01470_),
    .Z(_01471_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _05563_ (.A1(_01461_),
    .A2(\soc.spi_video_ram_1.buffer_index[1] ),
    .B(_01470_),
    .ZN(_01472_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _05564_ (.A1(_01468_),
    .A2(_01471_),
    .B(_01472_),
    .ZN(_01473_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05565_ (.I(\soc.spi_video_ram_1.buffer_index[5] ),
    .ZN(_01474_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _05566_ (.A1(_01460_),
    .A2(_01474_),
    .A3(_01464_),
    .ZN(_01475_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05567_ (.A1(\soc.spi_video_ram_1.buffer_index[1] ),
    .A2(_01475_),
    .ZN(_01476_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _05568_ (.A1(_01461_),
    .A2(_01476_),
    .ZN(_01477_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _05569_ (.A1(_01468_),
    .A2(\soc.spi_video_ram_1.output_buffer[12] ),
    .B1(_01477_),
    .B2(\soc.spi_video_ram_1.output_buffer[13] ),
    .ZN(_01478_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05570_ (.A1(_01467_),
    .A2(\soc.spi_video_ram_1.output_buffer[14] ),
    .ZN(_01479_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05571_ (.A1(\soc.spi_video_ram_1.output_buffer[15] ),
    .A2(_01475_),
    .ZN(_01480_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _05572_ (.A1(_01476_),
    .A2(_01479_),
    .B1(_01480_),
    .B2(_01467_),
    .ZN(_01481_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05573_ (.I(_01481_),
    .ZN(_01482_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _05574_ (.A1(_01467_),
    .A2(\soc.spi_video_ram_1.output_buffer[4] ),
    .B1(_01477_),
    .B2(\soc.spi_video_ram_1.output_buffer[5] ),
    .ZN(_01483_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _05575_ (.A1(_01468_),
    .A2(\soc.spi_video_ram_1.output_buffer[6] ),
    .B1(_01477_),
    .B2(\soc.spi_video_ram_1.output_buffer[7] ),
    .ZN(_01484_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _05576_ (.A1(_01461_),
    .A2(\soc.spi_video_ram_1.buffer_index[1] ),
    .Z(_01485_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _05577_ (.A1(_01462_),
    .A2(_01485_),
    .Z(_01486_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05578_ (.I(_01472_),
    .ZN(_01487_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _05579_ (.A1(_01463_),
    .A2(_01487_),
    .Z(_01488_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05580_ (.I0(_01478_),
    .I1(_01482_),
    .I2(_01483_),
    .I3(_01484_),
    .S0(_01486_),
    .S1(_01488_),
    .Z(_01489_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _05581_ (.I0(\soc.spi_video_ram_1.output_buffer[11] ),
    .I1(\soc.spi_video_ram_1.output_buffer[10] ),
    .S(_01461_),
    .Z(_01490_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _05582_ (.I0(\soc.spi_video_ram_1.output_buffer[9] ),
    .I1(\soc.spi_video_ram_1.output_buffer[8] ),
    .S(_01461_),
    .Z(_01491_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _05583_ (.A1(_01462_),
    .A2(_01485_),
    .ZN(_01492_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _05584_ (.I0(_01490_),
    .I1(_01491_),
    .S(_01492_),
    .Z(_01493_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05585_ (.A1(_01461_),
    .A2(\soc.spi_video_ram_1.buffer_index[1] ),
    .ZN(_01494_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _05586_ (.I0(\soc.spi_video_ram_1.output_buffer[3] ),
    .I1(\soc.spi_video_ram_1.output_buffer[2] ),
    .S(_01461_),
    .Z(_01495_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _05587_ (.A1(\soc.spi_video_ram_1.output_buffer[1] ),
    .A2(_01494_),
    .B1(_01486_),
    .B2(_01495_),
    .ZN(_01496_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05588_ (.A1(_01488_),
    .A2(_01496_),
    .ZN(_01497_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _05589_ (.A1(_01488_),
    .A2(_01493_),
    .B(_01473_),
    .C(_01497_),
    .ZN(_01498_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05590_ (.A1(_01473_),
    .A2(_01489_),
    .B(_01498_),
    .ZN(_01499_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _05591_ (.A1(_01460_),
    .A2(_01462_),
    .B(_01466_),
    .C(_01499_),
    .ZN(_01500_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05592_ (.I(_01467_),
    .Z(_01501_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _05593_ (.A1(_01501_),
    .A2(\soc.spi_video_ram_1.output_buffer[20] ),
    .B1(_01477_),
    .B2(\soc.spi_video_ram_1.output_buffer[21] ),
    .ZN(_01502_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _05594_ (.A1(_01501_),
    .A2(\soc.spi_video_ram_1.output_buffer[22] ),
    .B1(_01477_),
    .B2(\soc.spi_video_ram_1.output_buffer[23] ),
    .ZN(_01503_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05595_ (.A1(_01492_),
    .A2(_01503_),
    .ZN(_01504_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05596_ (.A1(_01473_),
    .A2(_01504_),
    .ZN(_01505_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05597_ (.A1(_01486_),
    .A2(_01502_),
    .B(_01505_),
    .ZN(_01506_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05598_ (.I(\soc.spi_video_ram_1.output_buffer[17] ),
    .ZN(_01507_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05599_ (.I(\soc.spi_video_ram_1.output_buffer[19] ),
    .ZN(_01508_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05600_ (.I(\soc.spi_video_ram_1.output_buffer[18] ),
    .ZN(_01509_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05601_ (.I(\soc.spi_video_ram_1.output_buffer[16] ),
    .ZN(_01510_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _05602_ (.I0(_01507_),
    .I1(_01508_),
    .I2(_01509_),
    .I3(_01510_),
    .S0(_01469_),
    .S1(_01501_),
    .Z(_01511_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05603_ (.A1(_01473_),
    .A2(_01511_),
    .ZN(_01512_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _05604_ (.A1(\soc.spi_video_ram_1.buffer_index[4] ),
    .A2(_01488_),
    .A3(_01506_),
    .A4(_01512_),
    .ZN(_01513_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05605_ (.A1(_01500_),
    .A2(_01513_),
    .ZN(_01514_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05606_ (.A1(_01428_),
    .A2(\soc.spi_video_ram_1.buffer_index[5] ),
    .ZN(_01515_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _05607_ (.A1(_01469_),
    .A2(_01470_),
    .ZN(_01516_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _05608_ (.I0(\soc.spi_video_ram_1.output_buffer[8] ),
    .I1(\soc.spi_video_ram_1.output_buffer[9] ),
    .S(_01468_),
    .Z(_01517_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05609_ (.I(_01470_),
    .ZN(_01518_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _05610_ (.A1(_01469_),
    .A2(_01518_),
    .Z(_01519_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _05611_ (.I0(\soc.spi_video_ram_1.output_buffer[10] ),
    .I1(\soc.spi_video_ram_1.output_buffer[11] ),
    .S(_01468_),
    .Z(_01520_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _05612_ (.A1(_01516_),
    .A2(_01517_),
    .B1(_01519_),
    .B2(_01520_),
    .ZN(_01521_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _05613_ (.I0(\soc.spi_video_ram_1.output_buffer[14] ),
    .I1(\soc.spi_video_ram_1.output_buffer[15] ),
    .S(_01468_),
    .Z(_01522_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _05614_ (.A1(_01469_),
    .A2(_01518_),
    .ZN(_01523_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _05615_ (.I0(\soc.spi_video_ram_1.output_buffer[12] ),
    .I1(\soc.spi_video_ram_1.output_buffer[13] ),
    .S(_01468_),
    .Z(_01524_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _05616_ (.A1(_01471_),
    .A2(_01522_),
    .B1(_01523_),
    .B2(_01524_),
    .ZN(_01525_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05617_ (.A1(_01521_),
    .A2(_01525_),
    .ZN(_01526_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05618_ (.A1(_01463_),
    .A2(_01526_),
    .ZN(_01527_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _05619_ (.I0(\soc.spi_video_ram_1.output_buffer[22] ),
    .I1(\soc.spi_video_ram_1.output_buffer[23] ),
    .S(_01468_),
    .Z(_01528_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05620_ (.A1(_01471_),
    .A2(_01528_),
    .ZN(_01529_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05621_ (.A1(_01467_),
    .A2(\soc.spi_video_ram_1.output_buffer[17] ),
    .ZN(_01530_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05622_ (.A1(_01468_),
    .A2(_01510_),
    .B(_01530_),
    .ZN(_01531_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05623_ (.A1(_01467_),
    .A2(\soc.spi_video_ram_1.output_buffer[18] ),
    .ZN(_01532_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05624_ (.A1(_01501_),
    .A2(_01508_),
    .B(_01532_),
    .ZN(_01533_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05625_ (.I(\soc.spi_video_ram_1.output_buffer[20] ),
    .ZN(_01534_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05626_ (.A1(_01467_),
    .A2(\soc.spi_video_ram_1.output_buffer[21] ),
    .ZN(_01535_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05627_ (.A1(_01501_),
    .A2(_01534_),
    .B(_01535_),
    .ZN(_01536_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _05628_ (.A1(_01516_),
    .A2(_01531_),
    .B1(_01533_),
    .B2(_01519_),
    .C1(_01523_),
    .C2(_01536_),
    .ZN(_01537_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _05629_ (.A1(\soc.spi_video_ram_1.buffer_index[4] ),
    .A2(_01529_),
    .A3(_01537_),
    .ZN(_01538_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05630_ (.I(\soc.spi_video_ram_1.output_buffer[4] ),
    .ZN(_01539_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05631_ (.A1(_01468_),
    .A2(\soc.spi_video_ram_1.output_buffer[5] ),
    .ZN(_01540_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _05632_ (.A1(_01501_),
    .A2(_01539_),
    .B(_01540_),
    .C(_01470_),
    .ZN(_01541_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05633_ (.I(_01541_),
    .ZN(_01542_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _05634_ (.A1(_01501_),
    .A2(\soc.spi_video_ram_1.output_buffer[1] ),
    .Z(_01543_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05635_ (.A1(_01470_),
    .A2(_01543_),
    .ZN(_01544_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _05636_ (.I0(\soc.spi_video_ram_1.output_buffer[2] ),
    .I1(\soc.spi_video_ram_1.output_buffer[3] ),
    .S(_01467_),
    .Z(_01545_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _05637_ (.I0(\soc.spi_video_ram_1.output_buffer[6] ),
    .I1(\soc.spi_video_ram_1.output_buffer[7] ),
    .S(_01467_),
    .Z(_01546_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _05638_ (.A1(_01519_),
    .A2(_01545_),
    .B1(_01546_),
    .B2(_01471_),
    .C(\soc.spi_video_ram_1.buffer_index[4] ),
    .ZN(_01547_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _05639_ (.A1(_01469_),
    .A2(_01542_),
    .A3(_01544_),
    .B(_01547_),
    .ZN(_01548_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05640_ (.A1(_01538_),
    .A2(_01548_),
    .ZN(_01549_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _05641_ (.A1(\soc.spi_video_ram_1.buffer_index[4] ),
    .A2(_01527_),
    .B1(_01549_),
    .B2(_01463_),
    .ZN(_01550_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _05642_ (.A1(_01514_),
    .A2(_01515_),
    .B1(_01550_),
    .B2(_01428_),
    .ZN(_01551_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05643_ (.I(_01551_),
    .ZN(net70));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _05644_ (.I(\soc.cpu.instruction[15] ),
    .Z(_01552_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05645_ (.I(_01552_),
    .Z(_01553_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05646_ (.I(\soc.cpu.DMuxJMP.sel[0] ),
    .ZN(_01554_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05647_ (.A1(_01552_),
    .A2(\soc.cpu.instruction[5] ),
    .ZN(_01555_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05648_ (.I(\soc.cpu.ALU.no ),
    .ZN(_01556_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _05649_ (.I(\soc.cpu.ALU.nx ),
    .Z(_01557_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _05650_ (.I(\soc.cpu.ALU.zx ),
    .ZN(_01558_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05651_ (.A1(_01558_),
    .A2(\soc.cpu.ALU.x[0] ),
    .ZN(_01559_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _05652_ (.A1(_01557_),
    .A2(_01559_),
    .Z(_01560_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05653_ (.I(\soc.cpu.ALU.ny ),
    .Z(_01561_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05654_ (.I(_01561_),
    .ZN(_01562_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _05655_ (.I(\soc.cpu.instruction[12] ),
    .ZN(_01563_));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 _05656_ (.I(\soc.cpu.AReg.data[0] ),
    .ZN(_01564_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05657_ (.I(\soc.cpu.AReg.data[1] ),
    .ZN(_01565_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05658_ (.A1(\soc.cpu.AReg.data[3] ),
    .A2(\soc.cpu.AReg.data[2] ),
    .ZN(_01566_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _05659_ (.A1(_01565_),
    .A2(_01566_),
    .ZN(_01567_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _05660_ (.A1(\soc.cpu.AReg.data[4] ),
    .A2(\soc.cpu.AReg.data[7] ),
    .A3(\soc.cpu.AReg.data[6] ),
    .ZN(_01568_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _05661_ (.A1(\soc.cpu.AReg.data[11] ),
    .A2(\soc.cpu.AReg.data[10] ),
    .A3(\soc.cpu.AReg.data[12] ),
    .A4(\soc.cpu.AReg.data[5] ),
    .ZN(_01569_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _05662_ (.A1(\soc.cpu.AReg.data[14] ),
    .A2(\soc.cpu.AReg.data[13] ),
    .Z(_01570_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05663_ (.A1(\soc.cpu.AReg.data[9] ),
    .A2(\soc.cpu.AReg.data[8] ),
    .ZN(_01571_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _05664_ (.A1(_01568_),
    .A2(_01569_),
    .A3(_01570_),
    .A4(_01571_),
    .ZN(_01572_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _05665_ (.A1(\soc.cpu.AReg.data[0] ),
    .A2(_01567_),
    .A3(_01572_),
    .ZN(_01573_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05666_ (.A1(net29),
    .A2(_01573_),
    .ZN(_01574_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _05667_ (.A1(_01564_),
    .A2(_01567_),
    .A3(_01572_),
    .ZN(_01575_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _05668_ (.A1(_01568_),
    .A2(_01569_),
    .A3(_01570_),
    .A4(_01571_),
    .Z(_01576_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _05669_ (.A1(\soc.cpu.AReg.data[1] ),
    .A2(_01566_),
    .Z(_01577_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _05670_ (.A1(net77),
    .A2(_01564_),
    .A3(_01576_),
    .A4(_01577_),
    .Z(_01578_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _05671_ (.A1(\soc.cpu.AReg.data[14] ),
    .A2(\soc.cpu.AReg.data[13] ),
    .ZN(_01579_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05672_ (.A1(\soc.ram_data_out[0] ),
    .A2(_01579_),
    .ZN(_01580_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05673_ (.A1(\soc.cpu.instruction[12] ),
    .A2(_01580_),
    .ZN(_01581_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _05674_ (.A1(\soc.gpio_i_stored[0] ),
    .A2(_01575_),
    .B(_01578_),
    .C(_01581_),
    .ZN(_01582_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _05675_ (.A1(_01563_),
    .A2(_01564_),
    .B1(_01574_),
    .B2(_01582_),
    .C(\soc.cpu.ALU.zy ),
    .ZN(_01583_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _05676_ (.A1(_01562_),
    .A2(_01583_),
    .Z(_01584_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05677_ (.I(\soc.cpu.ALU.f ),
    .Z(_01585_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _05678_ (.I(_01585_),
    .ZN(_01586_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05679_ (.A1(_01560_),
    .A2(_01584_),
    .B(_01586_),
    .ZN(_01587_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05680_ (.A1(_01560_),
    .A2(_01584_),
    .ZN(_01588_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _05681_ (.A1(_01556_),
    .A2(_01587_),
    .A3(_01588_),
    .Z(_01589_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05682_ (.I(\soc.cpu.instruction[5] ),
    .ZN(_01590_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _05683_ (.A1(\soc.cpu.instruction[15] ),
    .A2(_01590_),
    .ZN(_01591_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05684_ (.I(_01591_),
    .Z(_01592_));
 gf180mcu_fd_sc_mcu7t5v0__oai222_2 _05685_ (.A1(_01553_),
    .A2(_01554_),
    .B1(_01555_),
    .B2(_01589_),
    .C1(_01592_),
    .C2(_01564_),
    .ZN(\soc.cpu.PC.in[0] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _05686_ (.A1(\soc.cpu.instruction[15] ),
    .A2(\soc.cpu.instruction[5] ),
    .Z(_01593_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05687_ (.I(_01593_),
    .Z(_01594_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05688_ (.I(_01594_),
    .Z(_01595_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05689_ (.A1(_01558_),
    .A2(\soc.cpu.ALU.x[1] ),
    .ZN(_01596_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _05690_ (.A1(_01557_),
    .A2(_01596_),
    .Z(_01597_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05691_ (.I(\soc.cpu.instruction[12] ),
    .Z(_01598_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05692_ (.A1(\soc.ram_data_out[1] ),
    .A2(_01579_),
    .ZN(_01599_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05693_ (.A1(_01598_),
    .A2(_01599_),
    .ZN(_01600_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05694_ (.I(net38),
    .ZN(_01601_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _05695_ (.A1(net78),
    .A2(_01564_),
    .A3(_01576_),
    .A4(_01577_),
    .ZN(_01602_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _05696_ (.A1(\soc.cpu.AReg.data[3] ),
    .A2(\soc.cpu.AReg.data[2] ),
    .A3(\soc.cpu.AReg.data[1] ),
    .ZN(_01603_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _05697_ (.A1(\soc.gpio_i_stored[1] ),
    .A2(_01564_),
    .B(_01603_),
    .C(_01576_),
    .ZN(_01604_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _05698_ (.A1(_01601_),
    .A2(_01573_),
    .B1(_01602_),
    .B2(_01604_),
    .C(_01579_),
    .ZN(_01605_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _05699_ (.I(\soc.cpu.ALU.zy ),
    .ZN(_01606_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _05700_ (.A1(_01598_),
    .A2(\soc.cpu.AReg.data[1] ),
    .B1(_01600_),
    .B2(_01605_),
    .C(_01606_),
    .ZN(_01607_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _05701_ (.A1(_01561_),
    .A2(_01607_),
    .Z(_01608_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _05702_ (.A1(_01562_),
    .A2(_01597_),
    .A3(_01607_),
    .Z(_01609_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _05703_ (.A1(_01588_),
    .A2(_01609_),
    .ZN(_01610_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05704_ (.A1(_01585_),
    .A2(_01610_),
    .ZN(_01611_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _05705_ (.A1(_01585_),
    .A2(_01597_),
    .A3(_01608_),
    .B(_01611_),
    .ZN(_01612_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _05706_ (.A1(_01556_),
    .A2(_01612_),
    .Z(_01613_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _05707_ (.A1(_01553_),
    .A2(\soc.cpu.DMuxJMP.sel[1] ),
    .B1(\soc.cpu.AReg.data[1] ),
    .B2(_01592_),
    .ZN(_01614_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05708_ (.A1(_01595_),
    .A2(_01613_),
    .B(_01614_),
    .ZN(\soc.cpu.PC.in[1] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _05709_ (.I(\soc.cpu.ALU.no ),
    .Z(_01615_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05710_ (.A1(_01558_),
    .A2(\soc.cpu.ALU.x[2] ),
    .ZN(_01616_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _05711_ (.A1(_01557_),
    .A2(_01616_),
    .ZN(_01617_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05712_ (.I(_01563_),
    .Z(_01618_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05713_ (.I(\soc.cpu.AReg.data[2] ),
    .ZN(_01619_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05714_ (.A1(\soc.ram_data_out[2] ),
    .A2(_01579_),
    .B(_01563_),
    .ZN(_01620_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _05715_ (.A1(net79),
    .A2(_01564_),
    .A3(_01576_),
    .A4(_01577_),
    .Z(_01621_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _05716_ (.A1(\soc.gpio_i_stored[2] ),
    .A2(\soc.cpu.AReg.data[0] ),
    .A3(_01603_),
    .A4(_01576_),
    .Z(_01622_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _05717_ (.A1(\soc.cpu.AReg.data[0] ),
    .A2(net39),
    .A3(_01567_),
    .A4(_01572_),
    .Z(_01623_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _05718_ (.A1(_01573_),
    .A2(_01621_),
    .A3(_01622_),
    .B(_01623_),
    .ZN(_01624_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _05719_ (.A1(_01618_),
    .A2(_01619_),
    .B1(_01620_),
    .B2(_01624_),
    .C(\soc.cpu.ALU.zy ),
    .ZN(_01625_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _05720_ (.A1(_01561_),
    .A2(_01625_),
    .Z(_01626_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _05721_ (.A1(_01617_),
    .A2(_01626_),
    .Z(_01627_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _05722_ (.A1(_01560_),
    .A2(_01584_),
    .A3(_01609_),
    .B1(_01608_),
    .B2(_01597_),
    .ZN(_01628_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _05723_ (.A1(_01617_),
    .A2(_01626_),
    .A3(_01628_),
    .ZN(_01629_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05724_ (.A1(_01585_),
    .A2(_01629_),
    .ZN(_01630_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05725_ (.A1(_01585_),
    .A2(_01627_),
    .B(_01630_),
    .ZN(_01631_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _05726_ (.A1(_01615_),
    .A2(_01631_),
    .Z(_01632_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _05727_ (.A1(_01553_),
    .A2(\soc.cpu.DMuxJMP.sel[2] ),
    .B1(\soc.cpu.AReg.data[2] ),
    .B2(_01592_),
    .ZN(_01633_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05728_ (.A1(_01595_),
    .A2(_01632_),
    .B(_01633_),
    .ZN(\soc.cpu.PC.in[2] ));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _05729_ (.A1(_01617_),
    .A2(_01626_),
    .Z(_01634_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _05730_ (.A1(_01628_),
    .A2(_01634_),
    .B(_01627_),
    .ZN(_01635_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05731_ (.A1(_01558_),
    .A2(\soc.cpu.ALU.x[3] ),
    .ZN(_01636_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _05732_ (.A1(_01557_),
    .A2(_01636_),
    .ZN(_01637_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05733_ (.A1(\soc.ram_data_out[3] ),
    .A2(_01579_),
    .ZN(_01638_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05734_ (.A1(_01598_),
    .A2(_01638_),
    .ZN(_01639_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05735_ (.I(net40),
    .ZN(_01640_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05736_ (.A1(\soc.cpu.AReg.data[1] ),
    .A2(_01566_),
    .ZN(_01641_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _05737_ (.A1(\soc.cpu.AReg.data[0] ),
    .A2(_01572_),
    .A3(_01641_),
    .ZN(_01642_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _05738_ (.A1(net80),
    .A2(_01642_),
    .B1(_01575_),
    .B2(\soc.gpio_i_stored[3] ),
    .C(_01573_),
    .ZN(_01643_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05739_ (.A1(_01640_),
    .A2(_01573_),
    .B(_01643_),
    .ZN(_01644_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _05740_ (.A1(_01598_),
    .A2(\soc.cpu.AReg.data[3] ),
    .B1(_01639_),
    .B2(_01644_),
    .C(_01606_),
    .ZN(_01645_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _05741_ (.A1(_01562_),
    .A2(_01645_),
    .Z(_01646_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _05742_ (.A1(_01637_),
    .A2(_01646_),
    .ZN(_01647_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _05743_ (.A1(_01635_),
    .A2(_01647_),
    .Z(_01648_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05744_ (.A1(_01637_),
    .A2(_01646_),
    .ZN(_01649_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05745_ (.A1(_01586_),
    .A2(_01649_),
    .ZN(_01650_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05746_ (.A1(_01586_),
    .A2(_01648_),
    .B(_01650_),
    .ZN(_01651_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _05747_ (.A1(_01615_),
    .A2(_01651_),
    .Z(_01652_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _05748_ (.A1(_01553_),
    .A2(\soc.cpu.instruction[3] ),
    .B1(\soc.cpu.AReg.data[3] ),
    .B2(_01592_),
    .ZN(_01653_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05749_ (.A1(_01595_),
    .A2(_01652_),
    .B(_01653_),
    .ZN(\soc.cpu.PC.in[3] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _05750_ (.I(_01556_),
    .Z(_01654_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05751_ (.A1(_01558_),
    .A2(\soc.cpu.ALU.x[4] ),
    .ZN(_01655_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _05752_ (.A1(_01557_),
    .A2(_01655_),
    .ZN(_01656_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _05753_ (.A1(\soc.ram_data_out[4] ),
    .A2(_01579_),
    .B1(_01573_),
    .B2(net41),
    .C(_01563_),
    .ZN(_01657_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05754_ (.A1(_01598_),
    .A2(\soc.cpu.AReg.data[4] ),
    .B(_01606_),
    .ZN(_01658_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05755_ (.A1(_01657_),
    .A2(_01658_),
    .ZN(_01659_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _05756_ (.A1(_01561_),
    .A2(_01659_),
    .Z(_01660_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _05757_ (.A1(_01656_),
    .A2(_01660_),
    .Z(_01661_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _05758_ (.A1(_01635_),
    .A2(_01647_),
    .B(_01649_),
    .ZN(_01662_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _05759_ (.A1(_01656_),
    .A2(_01660_),
    .Z(_01663_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _05760_ (.A1(_01662_),
    .A2(_01663_),
    .Z(_01664_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _05761_ (.I0(_01661_),
    .I1(_01664_),
    .S(_01585_),
    .Z(_01665_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _05762_ (.A1(_01654_),
    .A2(_01665_),
    .Z(_01666_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _05763_ (.A1(_01553_),
    .A2(\soc.cpu.instruction[4] ),
    .B1(\soc.cpu.AReg.data[4] ),
    .B2(_01592_),
    .ZN(_01667_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05764_ (.A1(_01595_),
    .A2(_01666_),
    .B(_01667_),
    .ZN(\soc.cpu.PC.in[4] ));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _05765_ (.A1(_01662_),
    .A2(_01663_),
    .B(_01661_),
    .C(_01586_),
    .ZN(_01668_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05766_ (.I(_01585_),
    .Z(_01669_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05767_ (.I(_01558_),
    .Z(_01670_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05768_ (.A1(_01670_),
    .A2(\soc.cpu.ALU.x[5] ),
    .ZN(_01671_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _05769_ (.A1(_01557_),
    .A2(_01671_),
    .ZN(_01672_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _05770_ (.A1(\soc.ram_data_out[5] ),
    .A2(_01579_),
    .B1(_01573_),
    .B2(net42),
    .C(_01618_),
    .ZN(_01673_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05771_ (.A1(_01598_),
    .A2(\soc.cpu.AReg.data[5] ),
    .B(_01606_),
    .ZN(_01674_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05772_ (.A1(_01673_),
    .A2(_01674_),
    .ZN(_01675_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _05773_ (.A1(_01561_),
    .A2(_01675_),
    .Z(_01676_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05774_ (.A1(_01672_),
    .A2(_01676_),
    .ZN(_01677_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _05775_ (.A1(_01672_),
    .A2(_01676_),
    .Z(_01678_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05776_ (.A1(_01669_),
    .A2(_01677_),
    .B(_01678_),
    .ZN(_01679_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _05777_ (.A1(_01615_),
    .A2(_01668_),
    .A3(_01679_),
    .Z(_01680_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05778_ (.A1(_01553_),
    .A2(\soc.cpu.AReg.data[5] ),
    .ZN(_01681_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _05779_ (.A1(_01594_),
    .A2(_01680_),
    .B1(_01681_),
    .B2(_01590_),
    .ZN(\soc.cpu.PC.in[5] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05780_ (.I(_01586_),
    .Z(_01682_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05781_ (.A1(_01558_),
    .A2(\soc.cpu.ALU.x[6] ),
    .ZN(_01683_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _05782_ (.A1(_01557_),
    .A2(_01683_),
    .ZN(_01684_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _05783_ (.A1(\soc.ram_data_out[6] ),
    .A2(_01579_),
    .B1(_01573_),
    .B2(net43),
    .C(_01563_),
    .ZN(_01685_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05784_ (.A1(_01598_),
    .A2(\soc.cpu.AReg.data[6] ),
    .B(_01606_),
    .ZN(_01686_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05785_ (.A1(_01685_),
    .A2(_01686_),
    .ZN(_01687_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _05786_ (.A1(_01561_),
    .A2(_01687_),
    .Z(_01688_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _05787_ (.A1(_01684_),
    .A2(_01688_),
    .ZN(_01689_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05788_ (.A1(_01678_),
    .A2(_01677_),
    .ZN(_01690_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _05789_ (.A1(_01663_),
    .A2(_01690_),
    .Z(_01691_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _05790_ (.A1(_01656_),
    .A2(_01660_),
    .B1(_01672_),
    .B2(_01676_),
    .ZN(_01692_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05791_ (.A1(_01677_),
    .A2(_01692_),
    .ZN(_01693_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05792_ (.A1(_01662_),
    .A2(_01691_),
    .B(_01693_),
    .ZN(_01694_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _05793_ (.A1(_01689_),
    .A2(_01694_),
    .Z(_01695_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05794_ (.A1(_01684_),
    .A2(_01688_),
    .ZN(_01696_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05795_ (.A1(_01586_),
    .A2(_01696_),
    .ZN(_01697_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05796_ (.A1(_01682_),
    .A2(_01695_),
    .B(_01697_),
    .ZN(_01698_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _05797_ (.A1(_01615_),
    .A2(_01698_),
    .Z(_01699_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _05798_ (.A1(_01553_),
    .A2(_01615_),
    .B1(\soc.cpu.AReg.data[6] ),
    .B2(_01592_),
    .ZN(_01700_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05799_ (.A1(_01595_),
    .A2(_01699_),
    .B(_01700_),
    .ZN(\soc.cpu.PC.in[6] ));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _05800_ (.A1(_01689_),
    .A2(_01694_),
    .B(_01585_),
    .C(_01696_),
    .ZN(_01701_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _05801_ (.I(_01557_),
    .Z(_01702_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05802_ (.A1(_01670_),
    .A2(\soc.cpu.ALU.x[7] ),
    .ZN(_01703_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _05803_ (.A1(_01702_),
    .A2(_01703_),
    .ZN(_01704_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _05804_ (.I(_01561_),
    .Z(_01705_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _05805_ (.A1(\soc.ram_data_out[7] ),
    .A2(_01579_),
    .B1(_01573_),
    .B2(net44),
    .C(_01618_),
    .ZN(_01706_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05806_ (.A1(_01598_),
    .A2(\soc.cpu.AReg.data[7] ),
    .B(_01606_),
    .ZN(_01707_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05807_ (.A1(_01706_),
    .A2(_01707_),
    .ZN(_01708_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _05808_ (.A1(_01705_),
    .A2(_01708_),
    .Z(_01709_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05809_ (.A1(_01704_),
    .A2(_01709_),
    .ZN(_01710_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _05810_ (.A1(_01704_),
    .A2(_01709_),
    .Z(_01711_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05811_ (.A1(_01669_),
    .A2(_01710_),
    .B(_01711_),
    .ZN(_01712_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _05812_ (.A1(_01654_),
    .A2(_01701_),
    .A3(_01712_),
    .Z(_01713_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _05813_ (.A1(_01553_),
    .A2(_01669_),
    .B1(\soc.cpu.AReg.data[7] ),
    .B2(_01592_),
    .ZN(_01714_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05814_ (.A1(_01595_),
    .A2(_01713_),
    .B(_01714_),
    .ZN(\soc.cpu.PC.in[7] ));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05815_ (.A1(_01670_),
    .A2(\soc.cpu.ALU.x[8] ),
    .ZN(_01715_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _05816_ (.A1(_01702_),
    .A2(_01715_),
    .ZN(_01716_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05817_ (.I(\soc.cpu.ALU.zy ),
    .Z(_01717_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _05818_ (.A1(_01563_),
    .A2(_01570_),
    .ZN(_01718_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _05819_ (.A1(_01618_),
    .A2(\soc.cpu.AReg.data[8] ),
    .B1(_01718_),
    .B2(\soc.ram_data_out[8] ),
    .ZN(_01719_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05820_ (.A1(_01717_),
    .A2(_01719_),
    .ZN(_01720_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _05821_ (.A1(_01705_),
    .A2(_01720_),
    .Z(_01721_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05822_ (.A1(_01716_),
    .A2(_01721_),
    .ZN(_01722_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _05823_ (.A1(_01689_),
    .A2(_01711_),
    .A3(_01710_),
    .ZN(_01723_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _05824_ (.A1(_01662_),
    .A2(_01691_),
    .A3(_01723_),
    .ZN(_01724_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05825_ (.A1(_01693_),
    .A2(_01723_),
    .ZN(_01725_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05826_ (.A1(_01696_),
    .A2(_01710_),
    .ZN(_01726_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05827_ (.A1(_01711_),
    .A2(_01726_),
    .ZN(_01727_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _05828_ (.A1(_01725_),
    .A2(_01727_),
    .Z(_01728_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _05829_ (.A1(_01716_),
    .A2(_01721_),
    .Z(_01729_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05830_ (.I(_01729_),
    .ZN(_01730_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05831_ (.A1(_01724_),
    .A2(_01728_),
    .B(_01730_),
    .ZN(_01731_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _05832_ (.A1(_01662_),
    .A2(_01691_),
    .A3(_01723_),
    .Z(_01732_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05833_ (.A1(_01725_),
    .A2(_01727_),
    .ZN(_01733_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _05834_ (.A1(_01732_),
    .A2(_01733_),
    .A3(_01729_),
    .B(_01669_),
    .ZN(_01734_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _05835_ (.A1(_01669_),
    .A2(_01722_),
    .B1(_01731_),
    .B2(_01734_),
    .ZN(_01735_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _05836_ (.A1(_01654_),
    .A2(_01735_),
    .Z(_01736_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _05837_ (.A1(_01552_),
    .A2(_01705_),
    .B1(\soc.cpu.AReg.data[8] ),
    .B2(_01592_),
    .ZN(_01737_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05838_ (.A1(_01595_),
    .A2(_01736_),
    .B(_01737_),
    .ZN(\soc.cpu.PC.in[8] ));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05839_ (.A1(_01732_),
    .A2(_01733_),
    .B(_01729_),
    .ZN(_01738_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05840_ (.A1(_01670_),
    .A2(\soc.cpu.ALU.x[9] ),
    .ZN(_01739_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _05841_ (.A1(_01702_),
    .A2(_01739_),
    .ZN(_01740_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _05842_ (.A1(_01618_),
    .A2(\soc.cpu.AReg.data[9] ),
    .B1(_01718_),
    .B2(\soc.ram_data_out[9] ),
    .ZN(_01741_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05843_ (.A1(_01717_),
    .A2(_01741_),
    .ZN(_01742_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _05844_ (.A1(_01705_),
    .A2(_01742_),
    .Z(_01743_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05845_ (.A1(_01740_),
    .A2(_01743_),
    .ZN(_01744_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _05846_ (.A1(_01740_),
    .A2(_01743_),
    .Z(_01745_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _05847_ (.A1(_01744_),
    .A2(_01745_),
    .Z(_01746_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05848_ (.I(_01746_),
    .ZN(_01747_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05849_ (.A1(_01722_),
    .A2(_01738_),
    .B(_01747_),
    .ZN(_01748_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _05850_ (.A1(_01722_),
    .A2(_01738_),
    .A3(_01747_),
    .Z(_01749_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _05851_ (.A1(_01682_),
    .A2(_01740_),
    .A3(_01743_),
    .ZN(_01750_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _05852_ (.A1(_01682_),
    .A2(_01748_),
    .A3(_01749_),
    .B(_01750_),
    .ZN(_01751_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _05853_ (.A1(_01654_),
    .A2(_01751_),
    .Z(_01752_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _05854_ (.A1(_01552_),
    .A2(_01717_),
    .B1(\soc.cpu.AReg.data[9] ),
    .B2(_01592_),
    .ZN(_01753_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05855_ (.A1(_01595_),
    .A2(_01752_),
    .B(_01753_),
    .ZN(\soc.cpu.PC.in[9] ));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _05856_ (.A1(_01732_),
    .A2(_01733_),
    .B(_01729_),
    .C(_01746_),
    .ZN(_01754_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05857_ (.A1(_01722_),
    .A2(_01744_),
    .ZN(_01755_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05858_ (.A1(_01745_),
    .A2(_01755_),
    .ZN(_01756_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05859_ (.A1(_01670_),
    .A2(\soc.cpu.ALU.x[10] ),
    .ZN(_01757_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _05860_ (.A1(_01557_),
    .A2(_01757_),
    .ZN(_01758_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _05861_ (.A1(_01563_),
    .A2(\soc.cpu.AReg.data[10] ),
    .B1(_01718_),
    .B2(\soc.ram_data_out[10] ),
    .ZN(_01759_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05862_ (.A1(_01717_),
    .A2(_01759_),
    .ZN(_01760_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _05863_ (.A1(_01561_),
    .A2(_01760_),
    .Z(_01761_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _05864_ (.A1(_01758_),
    .A2(_01761_),
    .ZN(_01762_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05865_ (.A1(_01754_),
    .A2(_01756_),
    .B(_01762_),
    .ZN(_01763_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _05866_ (.A1(_01762_),
    .A2(_01754_),
    .A3(_01756_),
    .Z(_01764_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _05867_ (.A1(_01586_),
    .A2(_01758_),
    .A3(_01761_),
    .ZN(_01765_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _05868_ (.A1(_01682_),
    .A2(_01763_),
    .A3(_01764_),
    .B(_01765_),
    .ZN(_01766_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _05869_ (.A1(_01654_),
    .A2(_01766_),
    .Z(_01767_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _05870_ (.A1(_01552_),
    .A2(_01702_),
    .B1(\soc.cpu.AReg.data[10] ),
    .B2(_01591_),
    .ZN(_01768_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05871_ (.A1(_01595_),
    .A2(_01767_),
    .B(_01768_),
    .ZN(\soc.cpu.PC.in[10] ));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _05872_ (.A1(_01758_),
    .A2(_01761_),
    .B(_01763_),
    .C(_01682_),
    .ZN(_01769_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05873_ (.A1(_01670_),
    .A2(\soc.cpu.ALU.x[11] ),
    .ZN(_01770_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _05874_ (.A1(_01702_),
    .A2(_01770_),
    .ZN(_01771_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _05875_ (.A1(_01618_),
    .A2(\soc.cpu.AReg.data[11] ),
    .B1(_01718_),
    .B2(\soc.ram_data_out[11] ),
    .ZN(_01772_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05876_ (.A1(_01717_),
    .A2(_01772_),
    .ZN(_01773_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _05877_ (.A1(_01705_),
    .A2(_01773_),
    .Z(_01774_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05878_ (.A1(_01771_),
    .A2(_01774_),
    .ZN(_01775_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05879_ (.A1(_01771_),
    .A2(_01774_),
    .ZN(_01776_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05880_ (.A1(_01669_),
    .A2(_01776_),
    .ZN(_01777_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05881_ (.A1(_01775_),
    .A2(_01777_),
    .ZN(_01778_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _05882_ (.A1(_01654_),
    .A2(_01769_),
    .A3(_01778_),
    .Z(_01779_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _05883_ (.A1(_01552_),
    .A2(\soc.cpu.ALU.zx ),
    .B1(\soc.cpu.AReg.data[11] ),
    .B2(_01591_),
    .ZN(_01780_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05884_ (.A1(_01595_),
    .A2(_01779_),
    .B(_01780_),
    .ZN(\soc.cpu.PC.in[11] ));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05885_ (.A1(_01670_),
    .A2(\soc.cpu.ALU.x[12] ),
    .ZN(_01781_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _05886_ (.A1(_01702_),
    .A2(_01781_),
    .ZN(_01782_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _05887_ (.A1(_01618_),
    .A2(\soc.cpu.AReg.data[12] ),
    .B1(_01718_),
    .B2(\soc.ram_data_out[12] ),
    .ZN(_01783_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05888_ (.A1(_01717_),
    .A2(_01783_),
    .ZN(_01784_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _05889_ (.A1(_01705_),
    .A2(_01784_),
    .Z(_01785_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05890_ (.A1(_01782_),
    .A2(_01785_),
    .ZN(_01786_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05891_ (.A1(_01729_),
    .A2(_01746_),
    .ZN(_01787_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05892_ (.A1(_01762_),
    .A2(_01776_),
    .ZN(_01788_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05893_ (.A1(_01775_),
    .A2(_01788_),
    .ZN(_01789_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05894_ (.A1(_01787_),
    .A2(_01789_),
    .ZN(_01790_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05895_ (.A1(_01732_),
    .A2(_01733_),
    .B(_01790_),
    .ZN(_01791_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05896_ (.A1(_01758_),
    .A2(_01761_),
    .ZN(_01792_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05897_ (.A1(_01792_),
    .A2(_01776_),
    .B(_01775_),
    .ZN(_01793_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05898_ (.A1(_01756_),
    .A2(_01789_),
    .ZN(_01794_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05899_ (.A1(_01793_),
    .A2(_01794_),
    .ZN(_01795_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _05900_ (.A1(_01782_),
    .A2(_01785_),
    .Z(_01796_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05901_ (.I(_01796_),
    .ZN(_01797_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _05902_ (.A1(_01791_),
    .A2(_01795_),
    .B(_01797_),
    .ZN(_01798_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _05903_ (.A1(_01724_),
    .A2(_01728_),
    .B(_01787_),
    .C(_01789_),
    .ZN(_01799_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _05904_ (.A1(_01793_),
    .A2(_01794_),
    .Z(_01800_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _05905_ (.A1(_01799_),
    .A2(_01800_),
    .A3(_01796_),
    .B(_01669_),
    .ZN(_01801_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _05906_ (.A1(_01669_),
    .A2(_01786_),
    .B1(_01798_),
    .B2(_01801_),
    .ZN(_01802_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _05907_ (.A1(_01654_),
    .A2(_01802_),
    .Z(_01803_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _05908_ (.A1(_01552_),
    .A2(_01598_),
    .B1(\soc.cpu.AReg.data[12] ),
    .B2(_01591_),
    .ZN(_01804_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05909_ (.A1(_01594_),
    .A2(_01803_),
    .B(_01804_),
    .ZN(\soc.cpu.PC.in[12] ));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05910_ (.I(_01786_),
    .ZN(_01805_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05911_ (.A1(_01670_),
    .A2(\soc.cpu.ALU.x[13] ),
    .ZN(_01806_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _05912_ (.A1(_01702_),
    .A2(_01806_),
    .ZN(_01807_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _05913_ (.A1(_01618_),
    .A2(\soc.cpu.AReg.data[13] ),
    .B1(_01718_),
    .B2(\soc.ram_data_out[13] ),
    .ZN(_01808_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05914_ (.A1(_01717_),
    .A2(_01808_),
    .ZN(_01809_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _05915_ (.A1(_01705_),
    .A2(_01809_),
    .Z(_01810_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _05916_ (.A1(_01807_),
    .A2(_01810_),
    .Z(_01811_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _05917_ (.A1(_01805_),
    .A2(_01798_),
    .A3(_01811_),
    .ZN(_01812_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05918_ (.A1(_01799_),
    .A2(_01800_),
    .B(_01796_),
    .ZN(_01813_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05919_ (.I(_01811_),
    .ZN(_01814_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05920_ (.A1(_01786_),
    .A2(_01813_),
    .B(_01814_),
    .ZN(_01815_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _05921_ (.A1(_01807_),
    .A2(_01810_),
    .Z(_01816_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05922_ (.A1(_01682_),
    .A2(_01816_),
    .ZN(_01817_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _05923_ (.A1(_01682_),
    .A2(_01812_),
    .A3(_01815_),
    .B(_01817_),
    .ZN(_01818_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _05924_ (.A1(_01654_),
    .A2(_01818_),
    .Z(_01819_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _05925_ (.A1(_01552_),
    .A2(\soc.cpu.instruction[13] ),
    .B1(\soc.cpu.AReg.data[13] ),
    .B2(_01591_),
    .ZN(_01820_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05926_ (.A1(_01594_),
    .A2(_01819_),
    .B(_01820_),
    .ZN(\soc.cpu.PC.in[13] ));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05927_ (.A1(_01670_),
    .A2(\soc.cpu.ALU.x[14] ),
    .ZN(_01821_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _05928_ (.A1(_01702_),
    .A2(_01821_),
    .ZN(_01822_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _05929_ (.A1(_01618_),
    .A2(\soc.cpu.AReg.data[14] ),
    .B1(_01718_),
    .B2(\soc.ram_data_out[14] ),
    .ZN(_01823_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05930_ (.A1(_01717_),
    .A2(_01823_),
    .ZN(_01824_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _05931_ (.A1(_01705_),
    .A2(_01824_),
    .Z(_01825_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _05932_ (.A1(_01822_),
    .A2(_01825_),
    .Z(_01826_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _05933_ (.A1(_01816_),
    .A2(_01815_),
    .A3(_01826_),
    .ZN(_01827_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05934_ (.A1(_01807_),
    .A2(_01810_),
    .ZN(_01828_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05935_ (.A1(_01805_),
    .A2(_01798_),
    .B(_01811_),
    .ZN(_01829_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05936_ (.I(_01826_),
    .ZN(_01830_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05937_ (.A1(_01828_),
    .A2(_01829_),
    .B(_01830_),
    .ZN(_01831_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _05938_ (.A1(_01682_),
    .A2(_01822_),
    .A3(_01825_),
    .ZN(_01832_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _05939_ (.A1(_01682_),
    .A2(_01827_),
    .A3(_01831_),
    .B(_01832_),
    .ZN(_01833_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _05940_ (.A1(_01654_),
    .A2(_01833_),
    .Z(_01834_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _05941_ (.A1(_01552_),
    .A2(\soc.cpu.instruction[14] ),
    .B1(\soc.cpu.AReg.data[14] ),
    .B2(_01591_),
    .ZN(_01835_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05942_ (.A1(_01594_),
    .A2(_01834_),
    .B(_01835_),
    .ZN(\soc.cpu.PC.in[14] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05943_ (.I(\soc.video_generator_1.h_count[5] ),
    .Z(_01836_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _05944_ (.A1(\soc.video_generator_1.h_count[5] ),
    .A2(\soc.video_generator_1.h_count[6] ),
    .B(\soc.video_generator_1.h_count[7] ),
    .ZN(_01837_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _05945_ (.I(_01837_),
    .ZN(_01838_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _05946_ (.A1(\soc.video_generator_1.h_count[8] ),
    .A2(\soc.video_generator_1.h_count[9] ),
    .ZN(_01839_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _05947_ (.A1(_01838_),
    .A2(_01839_),
    .ZN(_01840_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _05948_ (.A1(_01836_),
    .A2(\soc.video_generator_1.h_count[7] ),
    .A3(\soc.video_generator_1.h_count[6] ),
    .B(_01840_),
    .ZN(_01841_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _05949_ (.A1(_01837_),
    .A2(_01839_),
    .ZN(_01842_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _05950_ (.A1(\soc.video_generator_1.h_count[3] ),
    .A2(\soc.video_generator_1.h_count[4] ),
    .A3(_01842_),
    .ZN(_01843_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _05951_ (.A1(\soc.video_generator_1.h_count[5] ),
    .A2(_01843_),
    .Z(_01844_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _05952_ (.A1(\soc.video_generator_1.h_count[5] ),
    .A2(\soc.video_generator_1.h_count[6] ),
    .ZN(_01845_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05953_ (.A1(_01842_),
    .A2(_01845_),
    .ZN(_01846_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _05954_ (.A1(_01844_),
    .A2(_01846_),
    .Z(_01847_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _05955_ (.A1(_01841_),
    .A2(_01847_),
    .Z(_01848_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _05956_ (.I(\soc.video_generator_1.v_count[6] ),
    .Z(_01849_));
 gf180mcu_fd_sc_mcu7t5v0__and4_4 _05957_ (.A1(\soc.video_generator_1.v_count[8] ),
    .A2(\soc.video_generator_1.v_count[7] ),
    .A3(_01849_),
    .A4(\soc.video_generator_1.v_count[5] ),
    .Z(_01850_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _05958_ (.A1(\soc.video_generator_1.v_count[2] ),
    .A2(\soc.video_generator_1.v_count[1] ),
    .Z(_01851_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _05959_ (.A1(\soc.video_generator_1.v_count[9] ),
    .A2(\soc.video_generator_1.v_count[3] ),
    .A3(_01850_),
    .A4(_01851_),
    .Z(_01852_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _05960_ (.I(\soc.video_generator_1.v_count[9] ),
    .Z(_01853_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _05961_ (.A1(\soc.video_generator_1.v_count[3] ),
    .A2(_01851_),
    .B(_01850_),
    .C(_01853_),
    .ZN(_01854_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _05962_ (.A1(_01852_),
    .A2(_01854_),
    .Z(_01855_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _05963_ (.A1(\soc.video_generator_1.v_count[7] ),
    .A2(_01849_),
    .A3(\soc.video_generator_1.v_count[5] ),
    .ZN(_01856_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _05964_ (.A1(\soc.video_generator_1.v_count[4] ),
    .A2(_01856_),
    .ZN(_01857_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05965_ (.A1(_01855_),
    .A2(_01857_),
    .ZN(_01858_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _05966_ (.A1(\soc.video_generator_1.v_count[9] ),
    .A2(_01850_),
    .A3(_01851_),
    .ZN(_01859_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_3 _05967_ (.I(\soc.video_generator_1.v_count[9] ),
    .ZN(_01860_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _05968_ (.I(\soc.video_generator_1.v_count[2] ),
    .ZN(_01861_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _05969_ (.I(\soc.video_generator_1.v_count[1] ),
    .ZN(_01862_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _05970_ (.A1(\soc.video_generator_1.v_count[8] ),
    .A2(\soc.video_generator_1.v_count[7] ),
    .A3(_01849_),
    .A4(\soc.video_generator_1.v_count[5] ),
    .ZN(_01863_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _05971_ (.A1(_01860_),
    .A2(_01861_),
    .A3(_01862_),
    .A4(_01863_),
    .ZN(_01864_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _05972_ (.A1(_01859_),
    .A2(_01864_),
    .Z(_01865_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _05973_ (.I(\soc.video_generator_1.v_count[0] ),
    .ZN(_01866_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _05974_ (.A1(_01860_),
    .A2(_01866_),
    .A3(_01863_),
    .A4(_01851_),
    .ZN(_01867_));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 _05975_ (.A1(_01852_),
    .A2(_01854_),
    .A3(_01857_),
    .A4(_01867_),
    .Z(_01868_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _05976_ (.A1(\soc.boot_loading_offset[1] ),
    .A2(_01860_),
    .A3(_01862_),
    .A4(_01863_),
    .ZN(_01869_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _05977_ (.A1(_01860_),
    .A2(_01866_),
    .A3(_01863_),
    .ZN(_01870_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05978_ (.I(\soc.boot_loading_offset[1] ),
    .ZN(_01871_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _05979_ (.A1(\soc.video_generator_1.v_count[9] ),
    .A2(\soc.video_generator_1.v_count[1] ),
    .A3(_01850_),
    .B(_01871_),
    .ZN(_01872_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _05980_ (.A1(\soc.boot_loading_offset[0] ),
    .A2(_01869_),
    .A3(_01870_),
    .A4(_01872_),
    .ZN(_01873_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05981_ (.A1(_01869_),
    .A2(_01873_),
    .ZN(_01874_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _05982_ (.A1(\soc.boot_loading_offset[2] ),
    .A2(_01865_),
    .A3(_01874_),
    .Z(_01875_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _05983_ (.A1(_01858_),
    .A2(_01865_),
    .B1(_01868_),
    .B2(_01875_),
    .ZN(_01876_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _05984_ (.A1(\soc.boot_loading_offset[2] ),
    .A2(_01859_),
    .A3(_01864_),
    .Z(_01877_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _05985_ (.A1(_01859_),
    .A2(_01864_),
    .B(\soc.boot_loading_offset[2] ),
    .ZN(_01878_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _05986_ (.A1(_01869_),
    .A2(_01873_),
    .B(_01878_),
    .ZN(_01879_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _05987_ (.A1(\soc.boot_loading_offset[3] ),
    .A2(_01877_),
    .A3(_01879_),
    .ZN(_01880_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05988_ (.I(\soc.boot_loading_offset[3] ),
    .ZN(_01881_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _05989_ (.A1(_01853_),
    .A2(\soc.video_generator_1.v_count[0] ),
    .A3(_01850_),
    .B(\soc.boot_loading_offset[0] ),
    .ZN(_01882_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05990_ (.I(_01882_),
    .ZN(_01883_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _05991_ (.A1(_01869_),
    .A2(_01872_),
    .Z(_01884_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _05992_ (.A1(\soc.video_generator_1.v_count[9] ),
    .A2(\soc.video_generator_1.v_count[1] ),
    .A3(_01850_),
    .ZN(_01885_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _05993_ (.A1(\soc.boot_loading_offset[1] ),
    .A2(_01885_),
    .Z(_01886_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _05994_ (.A1(_01883_),
    .A2(_01884_),
    .B(_01877_),
    .C(_01886_),
    .ZN(_01887_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _05995_ (.A1(_01881_),
    .A2(_01878_),
    .A3(_01887_),
    .B(_01868_),
    .ZN(_01888_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05996_ (.A1(_01880_),
    .A2(_01888_),
    .B(_01855_),
    .ZN(_01889_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _05997_ (.A1(_01876_),
    .A2(_01889_),
    .ZN(_01890_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _05998_ (.A1(\soc.video_generator_1.h_count[3] ),
    .A2(_01842_),
    .Z(_01891_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _05999_ (.A1(\soc.video_generator_1.h_count[3] ),
    .A2(\soc.video_generator_1.h_count[4] ),
    .B(_01842_),
    .ZN(_01892_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _06000_ (.A1(\soc.video_generator_1.h_count[4] ),
    .A2(_01891_),
    .B(_01892_),
    .ZN(_01893_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _06001_ (.A1(\soc.boot_loading_offset[0] ),
    .A2(_01870_),
    .A3(_01868_),
    .ZN(_01894_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06002_ (.I(\soc.boot_loading_offset[0] ),
    .ZN(_01895_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _06003_ (.A1(_01852_),
    .A2(_01854_),
    .A3(_01857_),
    .A4(_01867_),
    .ZN(_01896_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06004_ (.A1(_01860_),
    .A2(_01863_),
    .ZN(_01897_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06005_ (.A1(\soc.video_generator_1.v_count[0] ),
    .A2(_01897_),
    .ZN(_01898_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _06006_ (.A1(_01895_),
    .A2(_01896_),
    .B(_01898_),
    .ZN(_01899_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06007_ (.A1(_01893_),
    .A2(_01894_),
    .A3(_01899_),
    .ZN(_01900_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06008_ (.A1(\soc.video_generator_1.h_count[3] ),
    .A2(_01842_),
    .ZN(_01901_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _06009_ (.A1(\soc.display_clks_before_active[0] ),
    .A2(_01842_),
    .ZN(_01902_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06010_ (.A1(\soc.video_generator_1.h_count[1] ),
    .A2(_01842_),
    .ZN(_01903_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06011_ (.A1(\soc.video_generator_1.h_count[2] ),
    .A2(_01842_),
    .ZN(_01904_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _06012_ (.A1(_01902_),
    .A2(_01903_),
    .A3(_01904_),
    .ZN(_01905_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06013_ (.A1(_01901_),
    .A2(_01905_),
    .ZN(_01906_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _06014_ (.A1(_01894_),
    .A2(_01899_),
    .B(_01893_),
    .ZN(_01907_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _06015_ (.A1(_01900_),
    .A2(_01906_),
    .B(_01907_),
    .ZN(_01908_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06016_ (.A1(_01883_),
    .A2(_01884_),
    .Z(_01909_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06017_ (.A1(_01885_),
    .A2(_01858_),
    .B1(_01868_),
    .B2(_01909_),
    .ZN(_01910_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06018_ (.A1(_01837_),
    .A2(_01839_),
    .Z(_01911_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06019_ (.A1(_01836_),
    .A2(_01911_),
    .B(_01843_),
    .ZN(_01912_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06020_ (.A1(_01844_),
    .A2(_01912_),
    .ZN(_01913_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _06021_ (.A1(_01910_),
    .A2(_01913_),
    .ZN(_01914_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06022_ (.A1(_01910_),
    .A2(_01913_),
    .ZN(_01915_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _06023_ (.A1(_01908_),
    .A2(_01914_),
    .B(_01915_),
    .ZN(_01916_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _06024_ (.A1(_01844_),
    .A2(_01846_),
    .ZN(_01917_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06025_ (.A1(_01876_),
    .A2(_01917_),
    .Z(_01918_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06026_ (.A1(_01876_),
    .A2(_01917_),
    .ZN(_01919_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06027_ (.A1(_01916_),
    .A2(_01918_),
    .B(_01919_),
    .ZN(_01920_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _06028_ (.A1(_01848_),
    .A2(_01890_),
    .A3(_01920_),
    .Z(_01921_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06029_ (.A1(_01916_),
    .A2(_01918_),
    .Z(_01922_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _06030_ (.A1(_01908_),
    .A2(_01914_),
    .ZN(_01923_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06031_ (.I(_01923_),
    .Z(_01924_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06032_ (.A1(_01901_),
    .A2(_01905_),
    .Z(_01925_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06033_ (.I(\soc.video_generator_1.h_count[1] ),
    .ZN(_01926_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _06034_ (.A1(_01880_),
    .A2(_01888_),
    .B(_01855_),
    .C(_01876_),
    .ZN(_01927_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06035_ (.A1(_01881_),
    .A2(_01855_),
    .ZN(_01928_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _06036_ (.A1(_01881_),
    .A2(_01855_),
    .B1(_01878_),
    .B2(_01887_),
    .ZN(_01929_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _06037_ (.I(\soc.video_generator_1.v_count[4] ),
    .ZN(_01930_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _06038_ (.I(\soc.video_generator_1.v_count[3] ),
    .ZN(_01931_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _06039_ (.A1(_01930_),
    .A2(_01931_),
    .A3(_01859_),
    .ZN(_01932_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06040_ (.A1(\soc.video_generator_1.v_count[4] ),
    .A2(_01897_),
    .B(_01852_),
    .ZN(_01933_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06041_ (.A1(_01932_),
    .A2(_01933_),
    .Z(_01934_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _06042_ (.A1(\soc.boot_loading_offset[4] ),
    .A2(_01934_),
    .ZN(_01935_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _06043_ (.A1(_01928_),
    .A2(_01929_),
    .A3(_01935_),
    .Z(_01936_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06044_ (.A1(_01928_),
    .A2(_01929_),
    .B(_01935_),
    .ZN(_01937_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _06045_ (.A1(_01896_),
    .A2(_01936_),
    .A3(_01937_),
    .B(_01934_),
    .ZN(_01938_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06046_ (.I(\soc.video_generator_1.v_count[5] ),
    .Z(_01939_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06047_ (.A1(_01853_),
    .A2(_01850_),
    .ZN(_01940_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06048_ (.A1(_01939_),
    .A2(_01940_),
    .ZN(_01941_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06049_ (.A1(_01932_),
    .A2(_01941_),
    .Z(_01942_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _06050_ (.A1(_01868_),
    .A2(_01928_),
    .A3(_01929_),
    .A4(_01935_),
    .ZN(_01943_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06051_ (.A1(_01942_),
    .A2(_01943_),
    .ZN(_01944_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _06052_ (.A1(_01927_),
    .A2(_01938_),
    .B(_01944_),
    .ZN(_01945_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06053_ (.A1(_01927_),
    .A2(_01938_),
    .Z(_01946_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06054_ (.A1(_01841_),
    .A2(_01846_),
    .Z(_01947_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06055_ (.A1(\soc.video_generator_1.h_count[8] ),
    .A2(_01837_),
    .Z(_01948_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06056_ (.A1(\soc.video_generator_1.h_count[8] ),
    .A2(\soc.video_generator_1.h_count[9] ),
    .B(_01948_),
    .ZN(_01949_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06057_ (.A1(_01844_),
    .A2(_01947_),
    .B(_01949_),
    .ZN(_01950_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _06058_ (.A1(_01949_),
    .A2(_01844_),
    .A3(_01947_),
    .Z(_01951_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06059_ (.A1(_01950_),
    .A2(_01951_),
    .ZN(_01952_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06060_ (.A1(_01946_),
    .A2(_01952_),
    .ZN(_01953_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _06061_ (.A1(_01927_),
    .A2(_01938_),
    .A3(_01952_),
    .ZN(_01954_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06062_ (.A1(_01848_),
    .A2(_01890_),
    .ZN(_01955_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _06063_ (.A1(_01848_),
    .A2(_01890_),
    .B1(_01916_),
    .B2(_01918_),
    .C(_01919_),
    .ZN(_01956_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _06064_ (.A1(_01954_),
    .A2(_01955_),
    .A3(_01956_),
    .ZN(_01957_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _06065_ (.A1(_01927_),
    .A2(_01938_),
    .A3(_01944_),
    .Z(_01958_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _06066_ (.A1(\soc.video_generator_1.h_count[8] ),
    .A2(_01838_),
    .B(\soc.video_generator_1.h_count[9] ),
    .ZN(_01959_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06067_ (.A1(_01950_),
    .A2(_01959_),
    .Z(_01960_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _06068_ (.A1(_01945_),
    .A2(_01958_),
    .A3(_01960_),
    .ZN(_01961_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06069_ (.A1(_01945_),
    .A2(_01958_),
    .B(_01960_),
    .ZN(_01962_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _06070_ (.A1(_01953_),
    .A2(_01957_),
    .A3(_01961_),
    .B(_01962_),
    .ZN(_01963_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06071_ (.A1(_01853_),
    .A2(_01849_),
    .ZN(_01964_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06072_ (.A1(_01939_),
    .A2(_01940_),
    .A3(_01932_),
    .ZN(_01965_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06073_ (.I0(_01849_),
    .I1(_01964_),
    .S(_01965_),
    .Z(_01966_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _06074_ (.A1(_01945_),
    .A2(_01963_),
    .A3(_01966_),
    .Z(_01967_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06075_ (.A1(\soc.video_generator_1.h_count[1] ),
    .A2(\soc.display_clks_before_active[0] ),
    .ZN(_01968_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _06076_ (.A1(_01968_),
    .A2(_01904_),
    .B(_01905_),
    .ZN(_01969_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06077_ (.A1(_01891_),
    .A2(_01969_),
    .ZN(_01970_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _06078_ (.A1(_01926_),
    .A2(_01902_),
    .A3(_01967_),
    .A4(_01970_),
    .ZN(_01971_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06079_ (.A1(_01925_),
    .A2(_01971_),
    .ZN(_01972_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _06080_ (.A1(\soc.display_clks_before_active[0] ),
    .A2(\soc.video_generator_1.h_count[2] ),
    .A3(_01903_),
    .A4(_01967_),
    .Z(_01973_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06081_ (.A1(_01925_),
    .A2(_01973_),
    .Z(_01974_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _06082_ (.A1(_01893_),
    .A2(_01894_),
    .A3(_01899_),
    .Z(_01975_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06083_ (.A1(_01907_),
    .A2(_01975_),
    .ZN(_01976_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _06084_ (.A1(_01976_),
    .A2(_01906_),
    .Z(_01977_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06085_ (.A1(_01972_),
    .A2(_01974_),
    .B(_01977_),
    .ZN(_01978_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06086_ (.A1(_01924_),
    .A2(_01978_),
    .ZN(_01979_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06087_ (.A1(_01925_),
    .A2(_01969_),
    .B(_01970_),
    .ZN(_01980_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06088_ (.A1(_01967_),
    .A2(_01980_),
    .B(_01924_),
    .ZN(_01981_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _06089_ (.A1(\soc.video_generator_1.h_count[1] ),
    .A2(\soc.video_generator_1.h_count[2] ),
    .A3(_01901_),
    .ZN(_01982_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _06090_ (.A1(_01967_),
    .A2(_01982_),
    .Z(_01983_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06091_ (.A1(_01976_),
    .A2(_01983_),
    .ZN(_01984_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06092_ (.A1(_01977_),
    .A2(_01981_),
    .B(_01984_),
    .ZN(_01985_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _06093_ (.A1(_01891_),
    .A2(_01905_),
    .Z(_01986_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06094_ (.A1(_01902_),
    .A2(_01969_),
    .ZN(_01987_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06095_ (.I(_01987_),
    .ZN(_01988_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06096_ (.A1(_01902_),
    .A2(_01903_),
    .ZN(_01989_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06097_ (.A1(\soc.video_generator_1.h_count[1] ),
    .A2(\soc.display_clks_before_active[0] ),
    .ZN(_01990_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06098_ (.A1(_01989_),
    .A2(_01990_),
    .ZN(_01991_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06099_ (.A1(_01970_),
    .A2(_01991_),
    .ZN(_01992_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06100_ (.A1(\soc.video_generator_1.h_count[3] ),
    .A2(\soc.video_generator_1.h_count[2] ),
    .ZN(_01993_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06101_ (.I(\soc.display_clks_before_active[0] ),
    .ZN(_01994_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06102_ (.A1(\soc.display_clks_before_active[0] ),
    .A2(_01903_),
    .B(_01904_),
    .ZN(_01995_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06103_ (.A1(\soc.video_generator_1.h_count[1] ),
    .A2(_01994_),
    .B(_01995_),
    .ZN(_01996_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06104_ (.A1(_01989_),
    .A2(_01993_),
    .B1(_01996_),
    .B2(_01925_),
    .ZN(_01997_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06105_ (.I0(_01992_),
    .I1(_01997_),
    .S(_01923_),
    .Z(_01998_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _06106_ (.A1(_01902_),
    .A2(_01986_),
    .A3(_01924_),
    .B(_01998_),
    .ZN(_01999_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _06107_ (.A1(_01986_),
    .A2(_01988_),
    .B(_01999_),
    .C(_01967_),
    .ZN(_02000_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _06108_ (.A1(_01977_),
    .A2(_02000_),
    .B(_01978_),
    .C(_01922_),
    .ZN(_02001_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _06109_ (.A1(_01922_),
    .A2(_01979_),
    .A3(_01985_),
    .B(_02001_),
    .ZN(_02002_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _06110_ (.A1(_01921_),
    .A2(_02002_),
    .Z(_02003_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06111_ (.A1(_01924_),
    .A2(_01984_),
    .ZN(_02004_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06112_ (.A1(\soc.video_generator_1.h_count[2] ),
    .A2(_01902_),
    .ZN(_02005_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06113_ (.A1(_01926_),
    .A2(_02005_),
    .B(_01967_),
    .ZN(_02006_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06114_ (.A1(_01967_),
    .A2(_01988_),
    .B(_01986_),
    .ZN(_02007_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _06115_ (.A1(_01986_),
    .A2(_02006_),
    .B(_02007_),
    .C(_01977_),
    .ZN(_02008_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06116_ (.A1(_02004_),
    .A2(_02008_),
    .ZN(_02009_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _06117_ (.A1(_01907_),
    .A2(_01975_),
    .A3(_01983_),
    .B(_01924_),
    .ZN(_02010_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06118_ (.A1(_01922_),
    .A2(_02009_),
    .A3(_02010_),
    .ZN(_02011_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06119_ (.I(_01969_),
    .ZN(_02012_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06120_ (.A1(_01986_),
    .A2(_01924_),
    .B(_01991_),
    .ZN(_02013_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06121_ (.A1(_01976_),
    .A2(_01991_),
    .ZN(_02014_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06122_ (.A1(_02012_),
    .A2(_02013_),
    .B1(_02014_),
    .B2(_01925_),
    .ZN(_02015_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _06123_ (.A1(_01977_),
    .A2(_01924_),
    .A3(_01990_),
    .ZN(_02016_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06124_ (.A1(_01977_),
    .A2(_01924_),
    .ZN(_02017_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06125_ (.A1(_01977_),
    .A2(_01924_),
    .A3(_02005_),
    .ZN(_02018_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _06126_ (.A1(_01987_),
    .A2(_02017_),
    .B(_02018_),
    .C(_01989_),
    .ZN(_02019_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06127_ (.A1(_02016_),
    .A2(_02019_),
    .B(_01986_),
    .ZN(_02020_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06128_ (.A1(_01902_),
    .A2(_02015_),
    .B(_02020_),
    .ZN(_02021_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _06129_ (.A1(_01967_),
    .A2(_01922_),
    .A3(_02021_),
    .Z(_02022_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06130_ (.A1(_01921_),
    .A2(_02011_),
    .A3(_02022_),
    .ZN(_02023_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06131_ (.A1(_01955_),
    .A2(_01956_),
    .ZN(_02024_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _06132_ (.A1(_01954_),
    .A2(_02024_),
    .ZN(_02025_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06133_ (.A1(_02003_),
    .A2(_02023_),
    .B(_02025_),
    .ZN(_02026_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06134_ (.A1(_01953_),
    .A2(_01957_),
    .ZN(_02027_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _06135_ (.A1(_01945_),
    .A2(_01958_),
    .A3(_01960_),
    .Z(_02028_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06136_ (.A1(_02028_),
    .A2(_01962_),
    .Z(_02029_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06137_ (.A1(_01930_),
    .A2(_01931_),
    .B(_01940_),
    .ZN(_02030_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06138_ (.I(\soc.video_generator_1.h_count[7] ),
    .ZN(_02031_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _06139_ (.A1(_01891_),
    .A2(_01905_),
    .B(\soc.video_generator_1.h_count[4] ),
    .C(_02031_),
    .ZN(_02032_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _06140_ (.A1(_01836_),
    .A2(\soc.video_generator_1.h_count[6] ),
    .A3(_02032_),
    .Z(_02033_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06141_ (.I(\soc.video_generator_1.v_count[4] ),
    .Z(_02034_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06142_ (.A1(_02034_),
    .A2(\soc.video_generator_1.v_count[3] ),
    .A3(_01861_),
    .ZN(_02035_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _06143_ (.A1(\soc.video_generator_1.v_count[1] ),
    .A2(_01856_),
    .A3(_01897_),
    .A4(_02035_),
    .ZN(_02036_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06144_ (.A1(_01849_),
    .A2(_01939_),
    .A3(_01940_),
    .ZN(_02037_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06145_ (.A1(_01853_),
    .A2(\soc.video_generator_1.v_count[7] ),
    .B(_01959_),
    .ZN(_02038_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _06146_ (.A1(_01949_),
    .A2(_01893_),
    .A3(_02037_),
    .A4(_02038_),
    .Z(_02039_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _06147_ (.A1(_01870_),
    .A2(_02036_),
    .B(_02039_),
    .C(_01847_),
    .ZN(_02040_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _06148_ (.A1(_01947_),
    .A2(_02033_),
    .B(_02040_),
    .C(_01932_),
    .ZN(_02041_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _06149_ (.A1(_02027_),
    .A2(_02029_),
    .B1(_02030_),
    .B2(_01864_),
    .C(_02041_),
    .ZN(_02042_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06150_ (.A1(_01967_),
    .A2(_02005_),
    .ZN(_02043_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06151_ (.A1(_01977_),
    .A2(_02043_),
    .ZN(_02044_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06152_ (.A1(_01972_),
    .A2(_01973_),
    .B1(_02044_),
    .B2(_01925_),
    .ZN(_02045_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06153_ (.I(_01924_),
    .ZN(_02046_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06154_ (.A1(_01978_),
    .A2(_02045_),
    .B(_02046_),
    .ZN(_02047_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06155_ (.A1(_01922_),
    .A2(_02004_),
    .ZN(_02048_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06156_ (.A1(_01921_),
    .A2(_02048_),
    .ZN(_02049_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06157_ (.A1(_02047_),
    .A2(_02049_),
    .B(_02025_),
    .ZN(_02050_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _06158_ (.A1(_02027_),
    .A2(_02029_),
    .B(_02042_),
    .C(_02050_),
    .ZN(_02051_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _06159_ (.A1(_02026_),
    .A2(_02051_),
    .B(_01454_),
    .ZN(_02052_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _06160_ (.A1(\soc.hack_wait_clocks[1] ),
    .A2(\soc.hack_wait_clocks[0] ),
    .A3(_01452_),
    .A4(_01453_),
    .ZN(_02053_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06161_ (.A1(_01853_),
    .A2(\soc.video_generator_1.v_count[8] ),
    .ZN(_02054_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06162_ (.A1(_01853_),
    .A2(\soc.video_generator_1.v_count[7] ),
    .ZN(_02055_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _06163_ (.A1(_01849_),
    .A2(_01939_),
    .A3(_02034_),
    .A4(_01940_),
    .ZN(_02056_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06164_ (.A1(_02055_),
    .A2(_02056_),
    .Z(_02057_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06165_ (.A1(_02054_),
    .A2(_02057_),
    .Z(_02058_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06166_ (.A1(_01839_),
    .A2(_01846_),
    .ZN(_02059_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06167_ (.I0(\soc.spi_video_ram_1.read_value[2] ),
    .I1(\soc.spi_video_ram_1.read_value[3] ),
    .S(_01902_),
    .Z(_02060_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06168_ (.I(\soc.spi_video_ram_1.read_value[1] ),
    .ZN(_02061_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06169_ (.A1(_01994_),
    .A2(\soc.spi_video_ram_1.read_value[0] ),
    .ZN(_02062_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _06170_ (.A1(_02061_),
    .A2(_01902_),
    .B(_01903_),
    .C(_02062_),
    .ZN(_02063_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06171_ (.A1(_01949_),
    .A2(_01947_),
    .B1(_01959_),
    .B2(_01842_),
    .ZN(_02064_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _06172_ (.A1(_01903_),
    .A2(_02060_),
    .B(_02063_),
    .C(_02064_),
    .ZN(_02065_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _06173_ (.A1(_02053_),
    .A2(_02058_),
    .A3(_02059_),
    .A4(_02065_),
    .ZN(_02066_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _06174_ (.A1(_02052_),
    .A2(_02066_),
    .B(_01897_),
    .C(_01911_),
    .ZN(net76));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _06175_ (.I(\soc.ram_encoder_0.sram_sio_oe ),
    .ZN(net49));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _06176_ (.I(\soc.rom_encoder_0.sram_sio_oe ),
    .ZN(net53));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _06177_ (.I(\soc.spi_video_ram_1.sram_sio_oe ),
    .ZN(net57));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06178_ (.A1(\soc.video_generator_1.h_count[4] ),
    .A2(_01836_),
    .A3(\soc.video_generator_1.h_count[6] ),
    .ZN(_02067_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _06179_ (.A1(\soc.video_generator_1.h_count[4] ),
    .A2(_01836_),
    .A3(\soc.video_generator_1.h_count[6] ),
    .Z(_02068_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _06180_ (.A1(_02031_),
    .A2(_01839_),
    .A3(_02067_),
    .A4(_02068_),
    .ZN(net75));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06181_ (.A1(\soc.video_generator_1.v_count[8] ),
    .A2(\soc.video_generator_1.v_count[1] ),
    .ZN(_02069_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _06182_ (.A1(_01853_),
    .A2(_01931_),
    .A3(\soc.video_generator_1.v_count[2] ),
    .A4(_02069_),
    .ZN(_02070_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06183_ (.A1(_01857_),
    .A2(_02070_),
    .ZN(net74));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06184_ (.A1(_01516_),
    .A2(_01546_),
    .B(_01471_),
    .ZN(_02071_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _06185_ (.A1(_01469_),
    .A2(_01470_),
    .A3(_01463_),
    .ZN(_02072_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06186_ (.A1(_01460_),
    .A2(_02072_),
    .Z(_02073_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06187_ (.A1(_01463_),
    .A2(_01516_),
    .Z(_02074_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _06188_ (.A1(_01519_),
    .A2(_01543_),
    .B1(_01545_),
    .B2(_01523_),
    .C(_02074_),
    .ZN(_02075_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _06189_ (.A1(_01542_),
    .A2(_02071_),
    .B(_02073_),
    .C(_02075_),
    .ZN(_02076_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06190_ (.A1(_01471_),
    .A2(_01536_),
    .B1(_01531_),
    .B2(_01519_),
    .ZN(_02077_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06191_ (.A1(_01523_),
    .A2(_01533_),
    .B1(_01528_),
    .B2(_01516_),
    .ZN(_02078_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06192_ (.A1(_02077_),
    .A2(_02078_),
    .B(_02074_),
    .ZN(_02079_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _06193_ (.A1(_02073_),
    .A2(_02079_),
    .Z(_02080_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06194_ (.A1(_01516_),
    .A2(_01522_),
    .B1(_01524_),
    .B2(_01471_),
    .ZN(_02081_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _06195_ (.A1(_01476_),
    .A2(_02081_),
    .Z(_02082_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06196_ (.A1(_01520_),
    .A2(_01523_),
    .ZN(_02083_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06197_ (.A1(_01517_),
    .A2(_01519_),
    .ZN(_02084_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _06198_ (.A1(_02074_),
    .A2(_02082_),
    .A3(_02083_),
    .A4(_02084_),
    .ZN(_02085_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _06199_ (.A1(_01515_),
    .A2(_02076_),
    .A3(_02080_),
    .A4(_02085_),
    .Z(_02086_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06200_ (.I(_02086_),
    .Z(net71));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06201_ (.A1(_01470_),
    .A2(_01494_),
    .Z(_02087_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06202_ (.A1(_01492_),
    .A2(_01481_),
    .ZN(_02088_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _06203_ (.A1(_01492_),
    .A2(_01478_),
    .B(_02087_),
    .C(_02088_),
    .ZN(_02089_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06204_ (.A1(_01464_),
    .A2(_01494_),
    .ZN(_02090_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _06205_ (.A1(\soc.spi_video_ram_1.buffer_index[4] ),
    .A2(_02090_),
    .Z(_02091_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _06206_ (.A1(_01487_),
    .A2(_01490_),
    .B1(_01491_),
    .B2(_01486_),
    .C(_02087_),
    .ZN(_02092_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06207_ (.A1(_01470_),
    .A2(_01485_),
    .B(_01463_),
    .ZN(_02093_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06208_ (.A1(_02090_),
    .A2(_02093_),
    .Z(_02094_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06209_ (.A1(_02092_),
    .A2(_02094_),
    .ZN(_02095_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06210_ (.A1(_02089_),
    .A2(_02091_),
    .A3(_02095_),
    .ZN(_02096_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06211_ (.I0(\soc.spi_video_ram_1.output_buffer[19] ),
    .I1(\soc.spi_video_ram_1.output_buffer[16] ),
    .I2(\soc.spi_video_ram_1.output_buffer[17] ),
    .I3(\soc.spi_video_ram_1.output_buffer[18] ),
    .S0(_01501_),
    .S1(_01469_),
    .Z(_02097_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06212_ (.I(_02097_),
    .ZN(_02098_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06213_ (.A1(_01469_),
    .A2(\soc.spi_video_ram_1.output_buffer[1] ),
    .B(_01492_),
    .ZN(_02099_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06214_ (.A1(_01472_),
    .A2(_01495_),
    .B(_02091_),
    .ZN(_02100_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _06215_ (.A1(_02091_),
    .A2(_02098_),
    .B1(_02099_),
    .B2(_02100_),
    .ZN(_02101_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06216_ (.I0(_01502_),
    .I1(_01503_),
    .S(_01492_),
    .Z(_02102_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06217_ (.A1(_01486_),
    .A2(_01483_),
    .ZN(_02103_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06218_ (.A1(_01492_),
    .A2(_01484_),
    .ZN(_02104_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06219_ (.A1(_02091_),
    .A2(_02103_),
    .A3(_02104_),
    .ZN(_02105_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _06220_ (.A1(_02091_),
    .A2(_02102_),
    .B(_02105_),
    .C(_02087_),
    .ZN(_02106_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _06221_ (.A1(_02087_),
    .A2(_02101_),
    .B(_02106_),
    .C(_02094_),
    .ZN(_02107_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06222_ (.A1(\soc.spi_video_ram_1.buffer_index[4] ),
    .A2(_02090_),
    .B(\soc.spi_video_ram_1.buffer_index[5] ),
    .ZN(_02108_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06223_ (.A1(_01485_),
    .A2(_01475_),
    .B(_02108_),
    .ZN(_02109_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _06224_ (.A1(_02096_),
    .A2(_02107_),
    .B(_02109_),
    .C(_01428_),
    .ZN(net72));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _06225_ (.A1(_01428_),
    .A2(_01550_),
    .Z(_02110_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06226_ (.I(_02110_),
    .Z(net73));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _06227_ (.I(\soc.rom_encoder_0.toggled_sram_sck ),
    .ZN(_02111_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06228_ (.A1(net62),
    .A2(_02111_),
    .ZN(net63));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06229_ (.I(\soc.ram_encoder_0.toggled_sram_sck ),
    .ZN(_02112_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06230_ (.A1(net81),
    .A2(_02112_),
    .ZN(net82));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06231_ (.I(\soc.spi_video_ram_1.fifo_in_data[0] ),
    .Z(_02113_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06232_ (.A1(_01400_),
    .A2(_01405_),
    .ZN(_02114_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _06233_ (.I(\soc.spi_video_ram_1.write_fifo.write_pointer[4] ),
    .ZN(_02115_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06234_ (.I(\soc.spi_video_ram_1.write_fifo.write_pointer[2] ),
    .Z(_02116_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _06235_ (.A1(_02115_),
    .A2(_01403_),
    .A3(_02116_),
    .ZN(_02117_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06236_ (.A1(_02114_),
    .A2(_02117_),
    .ZN(_02118_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06237_ (.I(_02118_),
    .Z(_02119_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06238_ (.I(_02119_),
    .Z(_02120_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06239_ (.I0(_02113_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[18][0] ),
    .S(_02120_),
    .Z(_02121_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06240_ (.I(_02121_),
    .Z(_00012_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06241_ (.I(\soc.spi_video_ram_1.fifo_in_data[1] ),
    .Z(_02122_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06242_ (.I0(_02122_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[18][1] ),
    .S(_02120_),
    .Z(_02123_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06243_ (.I(_02123_),
    .Z(_00013_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06244_ (.I(\soc.spi_video_ram_1.fifo_in_data[2] ),
    .Z(_02124_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06245_ (.I0(_02124_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[18][2] ),
    .S(_02120_),
    .Z(_02125_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06246_ (.I(_02125_),
    .Z(_00014_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06247_ (.I(\soc.spi_video_ram_1.fifo_in_data[3] ),
    .Z(_02126_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06248_ (.I0(_02126_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[18][3] ),
    .S(_02120_),
    .Z(_02127_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06249_ (.I(_02127_),
    .Z(_00015_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06250_ (.I(\soc.spi_video_ram_1.fifo_in_data[4] ),
    .Z(_02128_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06251_ (.I0(_02128_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[18][4] ),
    .S(_02120_),
    .Z(_02129_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06252_ (.I(_02129_),
    .Z(_00016_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06253_ (.I(\soc.spi_video_ram_1.fifo_in_data[5] ),
    .Z(_02130_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06254_ (.I0(_02130_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[18][5] ),
    .S(_02120_),
    .Z(_02131_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06255_ (.I(_02131_),
    .Z(_00017_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06256_ (.I(\soc.spi_video_ram_1.fifo_in_data[6] ),
    .Z(_02132_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06257_ (.I0(_02132_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[18][6] ),
    .S(_02120_),
    .Z(_02133_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06258_ (.I(_02133_),
    .Z(_00018_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06259_ (.I(\soc.spi_video_ram_1.fifo_in_data[7] ),
    .Z(_02134_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06260_ (.I0(_02134_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[18][7] ),
    .S(_02120_),
    .Z(_02135_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06261_ (.I(_02135_),
    .Z(_00019_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06262_ (.I(\soc.spi_video_ram_1.fifo_in_data[8] ),
    .Z(_02136_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06263_ (.I0(_02136_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[18][8] ),
    .S(_02120_),
    .Z(_02137_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06264_ (.I(_02137_),
    .Z(_00020_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06265_ (.I(\soc.spi_video_ram_1.fifo_in_data[9] ),
    .Z(_02138_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06266_ (.I0(_02138_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[18][9] ),
    .S(_02120_),
    .Z(_02139_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06267_ (.I(_02139_),
    .Z(_00021_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06268_ (.I(\soc.spi_video_ram_1.fifo_in_data[10] ),
    .Z(_02140_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06269_ (.I(_02118_),
    .Z(_02141_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06270_ (.I0(_02140_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[18][10] ),
    .S(_02141_),
    .Z(_02142_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06271_ (.I(_02142_),
    .Z(_00022_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06272_ (.I(\soc.spi_video_ram_1.fifo_in_data[11] ),
    .Z(_02143_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06273_ (.I0(_02143_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[18][11] ),
    .S(_02141_),
    .Z(_02144_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06274_ (.I(_02144_),
    .Z(_00023_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06275_ (.I(\soc.spi_video_ram_1.fifo_in_data[12] ),
    .Z(_02145_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06276_ (.I0(_02145_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[18][12] ),
    .S(_02141_),
    .Z(_02146_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06277_ (.I(_02146_),
    .Z(_00024_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06278_ (.I(\soc.spi_video_ram_1.fifo_in_data[13] ),
    .Z(_02147_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06279_ (.I0(_02147_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[18][13] ),
    .S(_02141_),
    .Z(_02148_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06280_ (.I(_02148_),
    .Z(_00025_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06281_ (.I(\soc.spi_video_ram_1.fifo_in_data[14] ),
    .Z(_02149_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06282_ (.I0(_02149_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[18][14] ),
    .S(_02141_),
    .Z(_02150_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06283_ (.I(_02150_),
    .Z(_00026_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06284_ (.I(\soc.spi_video_ram_1.fifo_in_data[15] ),
    .Z(_02151_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06285_ (.I0(_02151_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[18][15] ),
    .S(_02141_),
    .Z(_02152_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06286_ (.I(_02152_),
    .Z(_00027_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06287_ (.I(\soc.spi_video_ram_1.fifo_in_address[0] ),
    .Z(_02153_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06288_ (.I0(_02153_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[18][16] ),
    .S(_02141_),
    .Z(_02154_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06289_ (.I(_02154_),
    .Z(_00028_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06290_ (.I(\soc.spi_video_ram_1.fifo_in_address[1] ),
    .Z(_02155_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06291_ (.I0(_02155_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[18][17] ),
    .S(_02141_),
    .Z(_02156_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06292_ (.I(_02156_),
    .Z(_00029_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06293_ (.I(\soc.spi_video_ram_1.fifo_in_address[2] ),
    .Z(_02157_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06294_ (.I0(_02157_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[18][18] ),
    .S(_02141_),
    .Z(_02158_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06295_ (.I(_02158_),
    .Z(_00030_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06296_ (.I(\soc.spi_video_ram_1.fifo_in_address[3] ),
    .Z(_02159_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06297_ (.I0(_02159_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[18][19] ),
    .S(_02141_),
    .Z(_02160_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06298_ (.I(_02160_),
    .Z(_00031_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06299_ (.I(\soc.spi_video_ram_1.fifo_in_address[4] ),
    .Z(_02161_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06300_ (.I0(_02161_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[18][20] ),
    .S(_02119_),
    .Z(_02162_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06301_ (.I(_02162_),
    .Z(_00032_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06302_ (.I(\soc.spi_video_ram_1.fifo_in_address[5] ),
    .Z(_02163_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06303_ (.I0(_02163_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[18][21] ),
    .S(_02119_),
    .Z(_02164_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06304_ (.I(_02164_),
    .Z(_00033_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06305_ (.I(\soc.spi_video_ram_1.fifo_in_address[6] ),
    .Z(_02165_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06306_ (.I0(_02165_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[18][22] ),
    .S(_02119_),
    .Z(_02166_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06307_ (.I(_02166_),
    .Z(_00034_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06308_ (.I(\soc.spi_video_ram_1.fifo_in_address[7] ),
    .Z(_02167_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06309_ (.I0(_02167_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[18][23] ),
    .S(_02119_),
    .Z(_02168_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06310_ (.I(_02168_),
    .Z(_00035_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06311_ (.I(\soc.spi_video_ram_1.fifo_in_address[8] ),
    .Z(_02169_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06312_ (.I0(_02169_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[18][24] ),
    .S(_02119_),
    .Z(_02170_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06313_ (.I(_02170_),
    .Z(_00036_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06314_ (.I(\soc.spi_video_ram_1.fifo_in_address[9] ),
    .Z(_02171_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06315_ (.I0(_02171_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[18][25] ),
    .S(_02119_),
    .Z(_02172_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06316_ (.I(_02172_),
    .Z(_00037_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06317_ (.I(\soc.spi_video_ram_1.fifo_in_address[10] ),
    .Z(_02173_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06318_ (.I0(_02173_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[18][26] ),
    .S(_02119_),
    .Z(_02174_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06319_ (.I(_02174_),
    .Z(_00038_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06320_ (.I(\soc.spi_video_ram_1.fifo_in_address[11] ),
    .Z(_02175_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06321_ (.I0(_02175_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[18][27] ),
    .S(_02119_),
    .Z(_02176_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06322_ (.I(_02176_),
    .Z(_00039_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06323_ (.I(\soc.spi_video_ram_1.fifo_in_address[12] ),
    .Z(_02177_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06324_ (.I0(_02177_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[18][28] ),
    .S(_02119_),
    .Z(_02178_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06325_ (.I(_02178_),
    .Z(_00040_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06326_ (.A1(\soc.spi_video_ram_1.write_fifo.write_pointer[1] ),
    .A2(_01444_),
    .ZN(_02179_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06327_ (.A1(_02117_),
    .A2(_02179_),
    .ZN(_02180_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06328_ (.I(_02180_),
    .Z(_02181_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06329_ (.I(_02181_),
    .Z(_02182_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06330_ (.I0(_02113_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[17][0] ),
    .S(_02182_),
    .Z(_02183_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06331_ (.I(_02183_),
    .Z(_00041_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06332_ (.I0(_02122_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[17][1] ),
    .S(_02182_),
    .Z(_02184_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06333_ (.I(_02184_),
    .Z(_00042_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06334_ (.I0(_02124_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[17][2] ),
    .S(_02182_),
    .Z(_02185_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06335_ (.I(_02185_),
    .Z(_00043_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06336_ (.I0(_02126_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[17][3] ),
    .S(_02182_),
    .Z(_02186_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06337_ (.I(_02186_),
    .Z(_00044_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06338_ (.I0(_02128_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[17][4] ),
    .S(_02182_),
    .Z(_02187_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06339_ (.I(_02187_),
    .Z(_00045_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06340_ (.I0(_02130_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[17][5] ),
    .S(_02182_),
    .Z(_02188_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06341_ (.I(_02188_),
    .Z(_00046_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06342_ (.I0(_02132_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[17][6] ),
    .S(_02182_),
    .Z(_02189_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06343_ (.I(_02189_),
    .Z(_00047_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06344_ (.I0(_02134_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[17][7] ),
    .S(_02182_),
    .Z(_02190_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06345_ (.I(_02190_),
    .Z(_00048_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06346_ (.I0(_02136_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[17][8] ),
    .S(_02182_),
    .Z(_02191_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06347_ (.I(_02191_),
    .Z(_00049_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06348_ (.I0(_02138_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[17][9] ),
    .S(_02182_),
    .Z(_02192_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06349_ (.I(_02192_),
    .Z(_00050_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06350_ (.I(_02180_),
    .Z(_02193_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06351_ (.I0(_02140_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[17][10] ),
    .S(_02193_),
    .Z(_02194_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06352_ (.I(_02194_),
    .Z(_00051_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06353_ (.I0(_02143_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[17][11] ),
    .S(_02193_),
    .Z(_02195_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06354_ (.I(_02195_),
    .Z(_00052_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06355_ (.I0(_02145_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[17][12] ),
    .S(_02193_),
    .Z(_02196_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06356_ (.I(_02196_),
    .Z(_00053_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06357_ (.I0(_02147_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[17][13] ),
    .S(_02193_),
    .Z(_02197_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06358_ (.I(_02197_),
    .Z(_00054_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06359_ (.I0(_02149_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[17][14] ),
    .S(_02193_),
    .Z(_02198_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06360_ (.I(_02198_),
    .Z(_00055_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06361_ (.I0(_02151_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[17][15] ),
    .S(_02193_),
    .Z(_02199_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06362_ (.I(_02199_),
    .Z(_00056_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06363_ (.I0(_02153_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[17][16] ),
    .S(_02193_),
    .Z(_02200_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06364_ (.I(_02200_),
    .Z(_00057_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06365_ (.I0(_02155_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[17][17] ),
    .S(_02193_),
    .Z(_02201_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06366_ (.I(_02201_),
    .Z(_00058_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06367_ (.I0(_02157_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[17][18] ),
    .S(_02193_),
    .Z(_02202_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06368_ (.I(_02202_),
    .Z(_00059_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06369_ (.I0(_02159_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[17][19] ),
    .S(_02193_),
    .Z(_02203_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06370_ (.I(_02203_),
    .Z(_00060_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06371_ (.I0(_02161_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[17][20] ),
    .S(_02181_),
    .Z(_02204_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06372_ (.I(_02204_),
    .Z(_00061_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06373_ (.I0(_02163_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[17][21] ),
    .S(_02181_),
    .Z(_02205_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06374_ (.I(_02205_),
    .Z(_00062_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06375_ (.I0(_02165_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[17][22] ),
    .S(_02181_),
    .Z(_02206_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06376_ (.I(_02206_),
    .Z(_00063_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06377_ (.I0(_02167_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[17][23] ),
    .S(_02181_),
    .Z(_02207_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06378_ (.I(_02207_),
    .Z(_00064_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06379_ (.I0(_02169_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[17][24] ),
    .S(_02181_),
    .Z(_02208_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06380_ (.I(_02208_),
    .Z(_00065_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06381_ (.I0(_02171_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[17][25] ),
    .S(_02181_),
    .Z(_02209_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06382_ (.I(_02209_),
    .Z(_00066_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06383_ (.I0(_02173_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[17][26] ),
    .S(_02181_),
    .Z(_02210_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06384_ (.I(_02210_),
    .Z(_00067_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06385_ (.I0(_02175_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[17][27] ),
    .S(_02181_),
    .Z(_02211_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06386_ (.I(_02211_),
    .Z(_00068_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06387_ (.I0(_02177_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[17][28] ),
    .S(_02181_),
    .Z(_02212_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06388_ (.I(_02212_),
    .Z(_00069_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06389_ (.I(\soc.spi_video_ram_1.fifo_in_data[0] ),
    .Z(_02213_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _06390_ (.A1(\soc.spi_video_ram_1.write_fifo.write_pointer[1] ),
    .A2(_01405_),
    .ZN(_02214_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06391_ (.A1(_02117_),
    .A2(_02214_),
    .Z(_02215_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06392_ (.I(_02215_),
    .Z(_02216_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06393_ (.I(_02216_),
    .Z(_02217_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06394_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[16][0] ),
    .I1(_02213_),
    .S(_02217_),
    .Z(_02218_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06395_ (.I(_02218_),
    .Z(_00070_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06396_ (.I(\soc.spi_video_ram_1.fifo_in_data[1] ),
    .Z(_02219_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06397_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[16][1] ),
    .I1(_02219_),
    .S(_02217_),
    .Z(_02220_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06398_ (.I(_02220_),
    .Z(_00071_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06399_ (.I(\soc.spi_video_ram_1.fifo_in_data[2] ),
    .Z(_02221_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06400_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[16][2] ),
    .I1(_02221_),
    .S(_02217_),
    .Z(_02222_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06401_ (.I(_02222_),
    .Z(_00072_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06402_ (.I(\soc.spi_video_ram_1.fifo_in_data[3] ),
    .Z(_02223_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06403_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[16][3] ),
    .I1(_02223_),
    .S(_02217_),
    .Z(_02224_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06404_ (.I(_02224_),
    .Z(_00073_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06405_ (.I(\soc.spi_video_ram_1.fifo_in_data[4] ),
    .Z(_02225_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06406_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[16][4] ),
    .I1(_02225_),
    .S(_02217_),
    .Z(_02226_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06407_ (.I(_02226_),
    .Z(_00074_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06408_ (.I(\soc.spi_video_ram_1.fifo_in_data[5] ),
    .Z(_02227_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06409_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[16][5] ),
    .I1(_02227_),
    .S(_02217_),
    .Z(_02228_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06410_ (.I(_02228_),
    .Z(_00075_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06411_ (.I(\soc.spi_video_ram_1.fifo_in_data[6] ),
    .Z(_02229_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06412_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[16][6] ),
    .I1(_02229_),
    .S(_02217_),
    .Z(_02230_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06413_ (.I(_02230_),
    .Z(_00076_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06414_ (.I(\soc.spi_video_ram_1.fifo_in_data[7] ),
    .Z(_02231_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06415_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[16][7] ),
    .I1(_02231_),
    .S(_02217_),
    .Z(_02232_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06416_ (.I(_02232_),
    .Z(_00077_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06417_ (.I(\soc.spi_video_ram_1.fifo_in_data[8] ),
    .Z(_02233_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06418_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[16][8] ),
    .I1(_02233_),
    .S(_02217_),
    .Z(_02234_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06419_ (.I(_02234_),
    .Z(_00078_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06420_ (.I(\soc.spi_video_ram_1.fifo_in_data[9] ),
    .Z(_02235_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06421_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[16][9] ),
    .I1(_02235_),
    .S(_02217_),
    .Z(_02236_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06422_ (.I(_02236_),
    .Z(_00079_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06423_ (.I(\soc.spi_video_ram_1.fifo_in_data[10] ),
    .Z(_02237_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06424_ (.I(_02215_),
    .Z(_02238_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06425_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[16][10] ),
    .I1(_02237_),
    .S(_02238_),
    .Z(_02239_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06426_ (.I(_02239_),
    .Z(_00080_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06427_ (.I(\soc.spi_video_ram_1.fifo_in_data[11] ),
    .Z(_02240_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06428_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[16][11] ),
    .I1(_02240_),
    .S(_02238_),
    .Z(_02241_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06429_ (.I(_02241_),
    .Z(_00081_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06430_ (.I(\soc.spi_video_ram_1.fifo_in_data[12] ),
    .Z(_02242_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06431_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[16][12] ),
    .I1(_02242_),
    .S(_02238_),
    .Z(_02243_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06432_ (.I(_02243_),
    .Z(_00082_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06433_ (.I(\soc.spi_video_ram_1.fifo_in_data[13] ),
    .Z(_02244_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06434_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[16][13] ),
    .I1(_02244_),
    .S(_02238_),
    .Z(_02245_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06435_ (.I(_02245_),
    .Z(_00083_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06436_ (.I(\soc.spi_video_ram_1.fifo_in_data[14] ),
    .Z(_02246_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06437_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[16][14] ),
    .I1(_02246_),
    .S(_02238_),
    .Z(_02247_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06438_ (.I(_02247_),
    .Z(_00084_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06439_ (.I(\soc.spi_video_ram_1.fifo_in_data[15] ),
    .Z(_02248_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06440_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[16][15] ),
    .I1(_02248_),
    .S(_02238_),
    .Z(_02249_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06441_ (.I(_02249_),
    .Z(_00085_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06442_ (.I(\soc.spi_video_ram_1.fifo_in_address[0] ),
    .Z(_02250_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06443_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[16][16] ),
    .I1(_02250_),
    .S(_02238_),
    .Z(_02251_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06444_ (.I(_02251_),
    .Z(_00086_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06445_ (.I(\soc.spi_video_ram_1.fifo_in_address[1] ),
    .Z(_02252_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06446_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[16][17] ),
    .I1(_02252_),
    .S(_02238_),
    .Z(_02253_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06447_ (.I(_02253_),
    .Z(_00087_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06448_ (.I(\soc.spi_video_ram_1.fifo_in_address[2] ),
    .Z(_02254_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06449_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[16][18] ),
    .I1(_02254_),
    .S(_02238_),
    .Z(_02255_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06450_ (.I(_02255_),
    .Z(_00088_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06451_ (.I(\soc.spi_video_ram_1.fifo_in_address[3] ),
    .Z(_02256_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06452_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[16][19] ),
    .I1(_02256_),
    .S(_02238_),
    .Z(_02257_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06453_ (.I(_02257_),
    .Z(_00089_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06454_ (.I(\soc.spi_video_ram_1.fifo_in_address[4] ),
    .Z(_02258_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06455_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[16][20] ),
    .I1(_02258_),
    .S(_02216_),
    .Z(_02259_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06456_ (.I(_02259_),
    .Z(_00090_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06457_ (.I(\soc.spi_video_ram_1.fifo_in_address[5] ),
    .Z(_02260_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06458_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[16][21] ),
    .I1(_02260_),
    .S(_02216_),
    .Z(_02261_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06459_ (.I(_02261_),
    .Z(_00091_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06460_ (.I(\soc.spi_video_ram_1.fifo_in_address[6] ),
    .Z(_02262_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06461_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[16][22] ),
    .I1(_02262_),
    .S(_02216_),
    .Z(_02263_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06462_ (.I(_02263_),
    .Z(_00092_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06463_ (.I(\soc.spi_video_ram_1.fifo_in_address[7] ),
    .Z(_02264_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06464_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[16][23] ),
    .I1(_02264_),
    .S(_02216_),
    .Z(_02265_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06465_ (.I(_02265_),
    .Z(_00093_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06466_ (.I(\soc.spi_video_ram_1.fifo_in_address[8] ),
    .Z(_02266_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06467_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[16][24] ),
    .I1(_02266_),
    .S(_02216_),
    .Z(_02267_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06468_ (.I(_02267_),
    .Z(_00094_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06469_ (.I(\soc.spi_video_ram_1.fifo_in_address[9] ),
    .Z(_02268_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06470_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[16][25] ),
    .I1(_02268_),
    .S(_02216_),
    .Z(_02269_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06471_ (.I(_02269_),
    .Z(_00095_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06472_ (.I(\soc.spi_video_ram_1.fifo_in_address[10] ),
    .Z(_02270_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06473_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[16][26] ),
    .I1(_02270_),
    .S(_02216_),
    .Z(_02271_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06474_ (.I(_02271_),
    .Z(_00096_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06475_ (.I(\soc.spi_video_ram_1.fifo_in_address[11] ),
    .Z(_02272_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06476_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[16][27] ),
    .I1(_02272_),
    .S(_02216_),
    .Z(_02273_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06477_ (.I(_02273_),
    .Z(_00097_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06478_ (.I(\soc.spi_video_ram_1.fifo_in_address[12] ),
    .Z(_02274_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06479_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[16][28] ),
    .I1(_02274_),
    .S(_02216_),
    .Z(_02275_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06480_ (.I(_02275_),
    .Z(_00098_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _06481_ (.A1(\soc.spi_video_ram_1.write_fifo.write_pointer[4] ),
    .A2(_01403_),
    .A3(_02116_),
    .ZN(_02276_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06482_ (.A1(_02214_),
    .A2(_02276_),
    .ZN(_02277_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06483_ (.I(_02277_),
    .Z(_02278_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06484_ (.I(_02278_),
    .Z(_02279_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06485_ (.I0(_02113_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[0][0] ),
    .S(_02279_),
    .Z(_02280_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06486_ (.I(_02280_),
    .Z(_00099_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06487_ (.I0(_02122_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[0][1] ),
    .S(_02279_),
    .Z(_02281_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06488_ (.I(_02281_),
    .Z(_00100_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06489_ (.I0(_02124_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[0][2] ),
    .S(_02279_),
    .Z(_02282_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06490_ (.I(_02282_),
    .Z(_00101_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06491_ (.I0(_02126_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[0][3] ),
    .S(_02279_),
    .Z(_02283_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06492_ (.I(_02283_),
    .Z(_00102_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06493_ (.I0(_02128_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[0][4] ),
    .S(_02279_),
    .Z(_02284_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06494_ (.I(_02284_),
    .Z(_00103_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06495_ (.I0(_02130_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[0][5] ),
    .S(_02279_),
    .Z(_02285_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06496_ (.I(_02285_),
    .Z(_00104_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06497_ (.I0(_02132_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[0][6] ),
    .S(_02279_),
    .Z(_02286_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06498_ (.I(_02286_),
    .Z(_00105_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06499_ (.I0(_02134_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[0][7] ),
    .S(_02279_),
    .Z(_02287_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06500_ (.I(_02287_),
    .Z(_00106_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06501_ (.I0(_02136_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[0][8] ),
    .S(_02279_),
    .Z(_02288_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06502_ (.I(_02288_),
    .Z(_00107_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06503_ (.I0(_02138_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[0][9] ),
    .S(_02279_),
    .Z(_02289_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06504_ (.I(_02289_),
    .Z(_00108_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06505_ (.I(_02277_),
    .Z(_02290_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06506_ (.I0(_02140_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[0][10] ),
    .S(_02290_),
    .Z(_02291_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06507_ (.I(_02291_),
    .Z(_00109_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06508_ (.I0(_02143_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[0][11] ),
    .S(_02290_),
    .Z(_02292_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06509_ (.I(_02292_),
    .Z(_00110_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06510_ (.I0(_02145_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[0][12] ),
    .S(_02290_),
    .Z(_02293_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06511_ (.I(_02293_),
    .Z(_00111_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06512_ (.I0(_02147_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[0][13] ),
    .S(_02290_),
    .Z(_02294_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06513_ (.I(_02294_),
    .Z(_00112_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06514_ (.I0(_02149_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[0][14] ),
    .S(_02290_),
    .Z(_02295_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06515_ (.I(_02295_),
    .Z(_00113_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06516_ (.I0(_02151_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[0][15] ),
    .S(_02290_),
    .Z(_02296_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06517_ (.I(_02296_),
    .Z(_00114_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06518_ (.I0(_02153_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[0][16] ),
    .S(_02290_),
    .Z(_02297_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06519_ (.I(_02297_),
    .Z(_00115_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06520_ (.I0(_02155_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[0][17] ),
    .S(_02290_),
    .Z(_02298_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06521_ (.I(_02298_),
    .Z(_00116_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06522_ (.I0(_02157_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[0][18] ),
    .S(_02290_),
    .Z(_02299_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06523_ (.I(_02299_),
    .Z(_00117_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06524_ (.I0(_02159_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[0][19] ),
    .S(_02290_),
    .Z(_02300_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06525_ (.I(_02300_),
    .Z(_00118_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06526_ (.I0(_02161_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[0][20] ),
    .S(_02278_),
    .Z(_02301_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06527_ (.I(_02301_),
    .Z(_00119_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06528_ (.I0(_02163_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[0][21] ),
    .S(_02278_),
    .Z(_02302_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06529_ (.I(_02302_),
    .Z(_00120_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06530_ (.I0(_02165_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[0][22] ),
    .S(_02278_),
    .Z(_02303_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06531_ (.I(_02303_),
    .Z(_00121_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06532_ (.I0(_02167_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[0][23] ),
    .S(_02278_),
    .Z(_02304_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06533_ (.I(_02304_),
    .Z(_00122_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06534_ (.I0(_02169_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[0][24] ),
    .S(_02278_),
    .Z(_02305_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06535_ (.I(_02305_),
    .Z(_00123_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06536_ (.I0(_02171_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[0][25] ),
    .S(_02278_),
    .Z(_02306_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06537_ (.I(_02306_),
    .Z(_00124_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06538_ (.I0(_02173_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[0][26] ),
    .S(_02278_),
    .Z(_02307_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06539_ (.I(_02307_),
    .Z(_00125_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06540_ (.I0(_02175_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[0][27] ),
    .S(_02278_),
    .Z(_02308_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06541_ (.I(_02308_),
    .Z(_00126_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06542_ (.I0(_02177_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[0][28] ),
    .S(_02278_),
    .Z(_02309_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06543_ (.I(_02309_),
    .Z(_00127_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06544_ (.I(\soc.spi_video_ram_1.fifo_in_data[0] ),
    .Z(_02310_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06545_ (.A1(_01400_),
    .A2(_01405_),
    .ZN(_02311_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06546_ (.I(_01403_),
    .ZN(_02312_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06547_ (.A1(\soc.spi_video_ram_1.write_fifo.write_pointer[4] ),
    .A2(_02312_),
    .ZN(_02313_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06548_ (.A1(_02116_),
    .A2(_02313_),
    .ZN(_02314_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06549_ (.A1(_02311_),
    .A2(_02314_),
    .ZN(_02315_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06550_ (.I(_02315_),
    .Z(_02316_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06551_ (.I(_02316_),
    .Z(_02317_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06552_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[13][0] ),
    .I1(_02310_),
    .S(_02317_),
    .Z(_02318_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06553_ (.I(_02318_),
    .Z(_00128_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06554_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[13][1] ),
    .I1(_02219_),
    .S(_02317_),
    .Z(_02319_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06555_ (.I(_02319_),
    .Z(_00129_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06556_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[13][2] ),
    .I1(_02221_),
    .S(_02317_),
    .Z(_02320_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06557_ (.I(_02320_),
    .Z(_00130_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06558_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[13][3] ),
    .I1(_02223_),
    .S(_02317_),
    .Z(_02321_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06559_ (.I(_02321_),
    .Z(_00131_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06560_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[13][4] ),
    .I1(_02225_),
    .S(_02317_),
    .Z(_02322_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06561_ (.I(_02322_),
    .Z(_00132_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06562_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[13][5] ),
    .I1(_02227_),
    .S(_02317_),
    .Z(_02323_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06563_ (.I(_02323_),
    .Z(_00133_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06564_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[13][6] ),
    .I1(_02229_),
    .S(_02317_),
    .Z(_02324_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06565_ (.I(_02324_),
    .Z(_00134_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06566_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[13][7] ),
    .I1(_02231_),
    .S(_02317_),
    .Z(_02325_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06567_ (.I(_02325_),
    .Z(_00135_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06568_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[13][8] ),
    .I1(_02233_),
    .S(_02317_),
    .Z(_02326_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06569_ (.I(_02326_),
    .Z(_00136_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06570_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[13][9] ),
    .I1(_02235_),
    .S(_02317_),
    .Z(_02327_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06571_ (.I(_02327_),
    .Z(_00137_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06572_ (.I(_02315_),
    .Z(_02328_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06573_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[13][10] ),
    .I1(_02237_),
    .S(_02328_),
    .Z(_02329_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06574_ (.I(_02329_),
    .Z(_00138_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06575_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[13][11] ),
    .I1(_02240_),
    .S(_02328_),
    .Z(_02330_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06576_ (.I(_02330_),
    .Z(_00139_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06577_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[13][12] ),
    .I1(_02242_),
    .S(_02328_),
    .Z(_02331_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06578_ (.I(_02331_),
    .Z(_00140_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06579_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[13][13] ),
    .I1(_02244_),
    .S(_02328_),
    .Z(_02332_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06580_ (.I(_02332_),
    .Z(_00141_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06581_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[13][14] ),
    .I1(_02246_),
    .S(_02328_),
    .Z(_02333_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06582_ (.I(_02333_),
    .Z(_00142_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06583_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[13][15] ),
    .I1(_02248_),
    .S(_02328_),
    .Z(_02334_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06584_ (.I(_02334_),
    .Z(_00143_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06585_ (.I(\soc.spi_video_ram_1.fifo_in_address[0] ),
    .Z(_02335_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06586_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[13][16] ),
    .I1(_02335_),
    .S(_02328_),
    .Z(_02336_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06587_ (.I(_02336_),
    .Z(_00144_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06588_ (.I(\soc.spi_video_ram_1.fifo_in_address[1] ),
    .Z(_02337_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06589_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[13][17] ),
    .I1(_02337_),
    .S(_02328_),
    .Z(_02338_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06590_ (.I(_02338_),
    .Z(_00145_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06591_ (.I(\soc.spi_video_ram_1.fifo_in_address[2] ),
    .Z(_02339_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06592_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[13][18] ),
    .I1(_02339_),
    .S(_02328_),
    .Z(_02340_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06593_ (.I(_02340_),
    .Z(_00146_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06594_ (.I(\soc.spi_video_ram_1.fifo_in_address[3] ),
    .Z(_02341_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06595_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[13][19] ),
    .I1(_02341_),
    .S(_02328_),
    .Z(_02342_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06596_ (.I(_02342_),
    .Z(_00147_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06597_ (.I(\soc.spi_video_ram_1.fifo_in_address[4] ),
    .Z(_02343_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06598_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[13][20] ),
    .I1(_02343_),
    .S(_02316_),
    .Z(_02344_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06599_ (.I(_02344_),
    .Z(_00148_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06600_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[13][21] ),
    .I1(_02260_),
    .S(_02316_),
    .Z(_02345_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06601_ (.I(_02345_),
    .Z(_00149_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06602_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[13][22] ),
    .I1(_02262_),
    .S(_02316_),
    .Z(_02346_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06603_ (.I(_02346_),
    .Z(_00150_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06604_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[13][23] ),
    .I1(_02264_),
    .S(_02316_),
    .Z(_02347_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06605_ (.I(_02347_),
    .Z(_00151_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06606_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[13][24] ),
    .I1(_02266_),
    .S(_02316_),
    .Z(_02348_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06607_ (.I(_02348_),
    .Z(_00152_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06608_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[13][25] ),
    .I1(_02268_),
    .S(_02316_),
    .Z(_02349_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06609_ (.I(_02349_),
    .Z(_00153_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06610_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[13][26] ),
    .I1(_02270_),
    .S(_02316_),
    .Z(_02350_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06611_ (.I(_02350_),
    .Z(_00154_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06612_ (.I(\soc.spi_video_ram_1.fifo_in_address[11] ),
    .Z(_02351_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06613_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[13][27] ),
    .I1(_02351_),
    .S(_02316_),
    .Z(_02352_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06614_ (.I(_02352_),
    .Z(_00155_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06615_ (.I(\soc.spi_video_ram_1.fifo_in_address[12] ),
    .Z(_02353_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06616_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[13][28] ),
    .I1(_02353_),
    .S(_02316_),
    .Z(_02354_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06617_ (.I(_02354_),
    .Z(_00156_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _06618_ (.A1(_02116_),
    .A2(_02214_),
    .A3(_02313_),
    .ZN(_02355_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06619_ (.I(_02355_),
    .Z(_02356_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06620_ (.I(_02356_),
    .Z(_02357_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06621_ (.I0(_02113_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[12][0] ),
    .S(_02357_),
    .Z(_02358_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06622_ (.I(_02358_),
    .Z(_00157_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06623_ (.I0(_02122_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[12][1] ),
    .S(_02357_),
    .Z(_02359_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06624_ (.I(_02359_),
    .Z(_00158_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06625_ (.I0(_02124_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[12][2] ),
    .S(_02357_),
    .Z(_02360_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06626_ (.I(_02360_),
    .Z(_00159_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06627_ (.I0(_02126_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[12][3] ),
    .S(_02357_),
    .Z(_02361_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06628_ (.I(_02361_),
    .Z(_00160_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06629_ (.I0(_02128_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[12][4] ),
    .S(_02357_),
    .Z(_02362_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06630_ (.I(_02362_),
    .Z(_00161_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06631_ (.I0(_02130_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[12][5] ),
    .S(_02357_),
    .Z(_02363_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06632_ (.I(_02363_),
    .Z(_00162_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06633_ (.I0(_02132_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[12][6] ),
    .S(_02357_),
    .Z(_02364_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06634_ (.I(_02364_),
    .Z(_00163_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06635_ (.I0(_02134_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[12][7] ),
    .S(_02357_),
    .Z(_02365_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06636_ (.I(_02365_),
    .Z(_00164_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06637_ (.I0(_02136_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[12][8] ),
    .S(_02357_),
    .Z(_02366_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06638_ (.I(_02366_),
    .Z(_00165_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06639_ (.I0(_02138_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[12][9] ),
    .S(_02357_),
    .Z(_02367_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06640_ (.I(_02367_),
    .Z(_00166_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06641_ (.I(_02355_),
    .Z(_02368_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06642_ (.I0(_02140_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[12][10] ),
    .S(_02368_),
    .Z(_02369_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06643_ (.I(_02369_),
    .Z(_00167_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06644_ (.I0(_02143_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[12][11] ),
    .S(_02368_),
    .Z(_02370_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06645_ (.I(_02370_),
    .Z(_00168_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06646_ (.I0(_02145_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[12][12] ),
    .S(_02368_),
    .Z(_02371_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06647_ (.I(_02371_),
    .Z(_00169_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06648_ (.I0(_02147_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[12][13] ),
    .S(_02368_),
    .Z(_02372_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06649_ (.I(_02372_),
    .Z(_00170_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06650_ (.I0(_02149_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[12][14] ),
    .S(_02368_),
    .Z(_02373_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06651_ (.I(_02373_),
    .Z(_00171_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06652_ (.I0(_02151_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[12][15] ),
    .S(_02368_),
    .Z(_02374_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06653_ (.I(_02374_),
    .Z(_00172_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06654_ (.I0(_02153_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[12][16] ),
    .S(_02368_),
    .Z(_02375_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06655_ (.I(_02375_),
    .Z(_00173_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06656_ (.I0(_02155_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[12][17] ),
    .S(_02368_),
    .Z(_02376_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06657_ (.I(_02376_),
    .Z(_00174_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06658_ (.I0(_02157_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[12][18] ),
    .S(_02368_),
    .Z(_02377_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06659_ (.I(_02377_),
    .Z(_00175_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06660_ (.I0(_02159_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[12][19] ),
    .S(_02368_),
    .Z(_02378_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06661_ (.I(_02378_),
    .Z(_00176_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06662_ (.I0(_02161_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[12][20] ),
    .S(_02356_),
    .Z(_02379_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06663_ (.I(_02379_),
    .Z(_00177_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06664_ (.I0(_02163_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[12][21] ),
    .S(_02356_),
    .Z(_02380_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06665_ (.I(_02380_),
    .Z(_00178_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06666_ (.I0(_02165_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[12][22] ),
    .S(_02356_),
    .Z(_02381_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06667_ (.I(_02381_),
    .Z(_00179_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06668_ (.I0(_02167_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[12][23] ),
    .S(_02356_),
    .Z(_02382_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06669_ (.I(_02382_),
    .Z(_00180_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06670_ (.I0(_02169_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[12][24] ),
    .S(_02356_),
    .Z(_02383_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06671_ (.I(_02383_),
    .Z(_00181_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06672_ (.I0(_02171_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[12][25] ),
    .S(_02356_),
    .Z(_02384_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06673_ (.I(_02384_),
    .Z(_00182_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06674_ (.I0(_02173_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[12][26] ),
    .S(_02356_),
    .Z(_02385_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06675_ (.I(_02385_),
    .Z(_00183_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06676_ (.I0(_02175_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[12][27] ),
    .S(_02356_),
    .Z(_02386_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06677_ (.I(_02386_),
    .Z(_00184_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06678_ (.I0(_02177_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[12][28] ),
    .S(_02356_),
    .Z(_02387_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06679_ (.I(_02387_),
    .Z(_00185_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06680_ (.A1(\soc.spi_video_ram_1.write_fifo.write_pointer[1] ),
    .A2(_01444_),
    .ZN(_02388_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06681_ (.A1(_02388_),
    .A2(_02314_),
    .ZN(_02389_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06682_ (.I(_02389_),
    .Z(_02390_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06683_ (.I(_02390_),
    .Z(_02391_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06684_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[14][0] ),
    .I1(_02310_),
    .S(_02391_),
    .Z(_02392_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06685_ (.I(_02392_),
    .Z(_00186_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06686_ (.I(\soc.spi_video_ram_1.fifo_in_data[1] ),
    .Z(_02393_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06687_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[14][1] ),
    .I1(_02393_),
    .S(_02391_),
    .Z(_02394_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06688_ (.I(_02394_),
    .Z(_00187_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06689_ (.I(\soc.spi_video_ram_1.fifo_in_data[2] ),
    .Z(_02395_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06690_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[14][2] ),
    .I1(_02395_),
    .S(_02391_),
    .Z(_02396_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06691_ (.I(_02396_),
    .Z(_00188_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06692_ (.I(\soc.spi_video_ram_1.fifo_in_data[3] ),
    .Z(_02397_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06693_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[14][3] ),
    .I1(_02397_),
    .S(_02391_),
    .Z(_02398_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06694_ (.I(_02398_),
    .Z(_00189_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06695_ (.I(\soc.spi_video_ram_1.fifo_in_data[4] ),
    .Z(_02399_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06696_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[14][4] ),
    .I1(_02399_),
    .S(_02391_),
    .Z(_02400_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06697_ (.I(_02400_),
    .Z(_00190_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06698_ (.I(\soc.spi_video_ram_1.fifo_in_data[5] ),
    .Z(_02401_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06699_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[14][5] ),
    .I1(_02401_),
    .S(_02391_),
    .Z(_02402_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06700_ (.I(_02402_),
    .Z(_00191_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06701_ (.I(\soc.spi_video_ram_1.fifo_in_data[6] ),
    .Z(_02403_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06702_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[14][6] ),
    .I1(_02403_),
    .S(_02391_),
    .Z(_02404_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06703_ (.I(_02404_),
    .Z(_00192_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06704_ (.I(\soc.spi_video_ram_1.fifo_in_data[7] ),
    .Z(_02405_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06705_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[14][7] ),
    .I1(_02405_),
    .S(_02391_),
    .Z(_02406_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06706_ (.I(_02406_),
    .Z(_00193_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06707_ (.I(\soc.spi_video_ram_1.fifo_in_data[8] ),
    .Z(_02407_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06708_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[14][8] ),
    .I1(_02407_),
    .S(_02391_),
    .Z(_02408_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06709_ (.I(_02408_),
    .Z(_00194_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06710_ (.I(\soc.spi_video_ram_1.fifo_in_data[9] ),
    .Z(_02409_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06711_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[14][9] ),
    .I1(_02409_),
    .S(_02391_),
    .Z(_02410_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06712_ (.I(_02410_),
    .Z(_00195_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06713_ (.I(\soc.spi_video_ram_1.fifo_in_data[10] ),
    .Z(_02411_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06714_ (.I(_02389_),
    .Z(_02412_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06715_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[14][10] ),
    .I1(_02411_),
    .S(_02412_),
    .Z(_02413_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06716_ (.I(_02413_),
    .Z(_00196_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06717_ (.I(\soc.spi_video_ram_1.fifo_in_data[11] ),
    .Z(_02414_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06718_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[14][11] ),
    .I1(_02414_),
    .S(_02412_),
    .Z(_02415_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06719_ (.I(_02415_),
    .Z(_00197_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06720_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[14][12] ),
    .I1(_02242_),
    .S(_02412_),
    .Z(_02416_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06721_ (.I(_02416_),
    .Z(_00198_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06722_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[14][13] ),
    .I1(_02244_),
    .S(_02412_),
    .Z(_02417_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06723_ (.I(_02417_),
    .Z(_00199_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06724_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[14][14] ),
    .I1(_02246_),
    .S(_02412_),
    .Z(_02418_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06725_ (.I(_02418_),
    .Z(_00200_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06726_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[14][15] ),
    .I1(_02248_),
    .S(_02412_),
    .Z(_02419_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06727_ (.I(_02419_),
    .Z(_00201_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06728_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[14][16] ),
    .I1(_02335_),
    .S(_02412_),
    .Z(_02420_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06729_ (.I(_02420_),
    .Z(_00202_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06730_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[14][17] ),
    .I1(_02337_),
    .S(_02412_),
    .Z(_02421_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06731_ (.I(_02421_),
    .Z(_00203_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06732_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[14][18] ),
    .I1(_02339_),
    .S(_02412_),
    .Z(_02422_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06733_ (.I(_02422_),
    .Z(_00204_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06734_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[14][19] ),
    .I1(_02341_),
    .S(_02412_),
    .Z(_02423_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06735_ (.I(_02423_),
    .Z(_00205_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06736_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[14][20] ),
    .I1(_02343_),
    .S(_02390_),
    .Z(_02424_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06737_ (.I(_02424_),
    .Z(_00206_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06738_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[14][21] ),
    .I1(_02260_),
    .S(_02390_),
    .Z(_02425_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06739_ (.I(_02425_),
    .Z(_00207_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06740_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[14][22] ),
    .I1(_02262_),
    .S(_02390_),
    .Z(_02426_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06741_ (.I(_02426_),
    .Z(_00208_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06742_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[14][23] ),
    .I1(_02264_),
    .S(_02390_),
    .Z(_02427_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06743_ (.I(_02427_),
    .Z(_00209_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06744_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[14][24] ),
    .I1(_02266_),
    .S(_02390_),
    .Z(_02428_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06745_ (.I(_02428_),
    .Z(_00210_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06746_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[14][25] ),
    .I1(_02268_),
    .S(_02390_),
    .Z(_02429_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06747_ (.I(_02429_),
    .Z(_00211_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06748_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[14][26] ),
    .I1(_02270_),
    .S(_02390_),
    .Z(_02430_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06749_ (.I(_02430_),
    .Z(_00212_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06750_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[14][27] ),
    .I1(_02351_),
    .S(_02390_),
    .Z(_02431_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06751_ (.I(_02431_),
    .Z(_00213_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06752_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[14][28] ),
    .I1(_02353_),
    .S(_02390_),
    .Z(_02432_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06753_ (.I(_02432_),
    .Z(_00214_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 _06754_ (.I(\soc.rom_encoder_0.current_state[0] ),
    .Z(_02433_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_4 _06755_ (.I(\soc.rom_encoder_0.current_state[2] ),
    .ZN(_02434_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 _06756_ (.I(\soc.rom_encoder_0.current_state[1] ),
    .Z(_02435_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _06757_ (.I(_02435_),
    .ZN(_02436_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06758_ (.A1(_02434_),
    .A2(_02436_),
    .ZN(_02437_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06759_ (.A1(_02433_),
    .A2(_02437_),
    .Z(_02438_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06760_ (.I(\soc.rom_encoder_0.output_bits_left[3] ),
    .ZN(_02439_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06761_ (.A1(_02439_),
    .A2(\soc.rom_encoder_0.output_bits_left[2] ),
    .ZN(_02440_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _06762_ (.A1(\soc.rom_encoder_0.output_bits_left[4] ),
    .A2(_02440_),
    .ZN(_02441_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _06763_ (.A1(\soc.rom_encoder_0.current_state[2] ),
    .A2(_02436_),
    .ZN(_02442_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _06764_ (.A1(_02433_),
    .A2(_02442_),
    .ZN(_02443_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06765_ (.A1(_02434_),
    .A2(_02435_),
    .ZN(_02444_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _06766_ (.A1(_02433_),
    .A2(_02444_),
    .ZN(_02445_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _06767_ (.A1(\soc.rom_encoder_0.request_write ),
    .A2(_02443_),
    .B(_02445_),
    .ZN(_02446_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06768_ (.A1(_02435_),
    .A2(_02433_),
    .ZN(_02447_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _06769_ (.A1(_02441_),
    .A2(_02446_),
    .B(_02447_),
    .C(_02111_),
    .ZN(_02448_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _06770_ (.A1(\soc.rom_encoder_0.initializing_step[4] ),
    .A2(\soc.rom_encoder_0.initializing_step[3] ),
    .A3(\soc.rom_encoder_0.initializing_step[2] ),
    .A4(\soc.rom_encoder_0.initializing_step[1] ),
    .ZN(_02449_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06771_ (.A1(_02433_),
    .A2(_02449_),
    .ZN(_02450_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06772_ (.A1(_02437_),
    .A2(_02450_),
    .ZN(_02451_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06773_ (.A1(_02448_),
    .A2(_02451_),
    .ZN(_02452_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _06774_ (.A1(_02438_),
    .A2(_02452_),
    .Z(_02453_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06775_ (.I(_02433_),
    .Z(_02454_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _06776_ (.A1(_02434_),
    .A2(_02454_),
    .B1(_02442_),
    .B2(_02441_),
    .ZN(_02455_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06777_ (.A1(\soc.rom_encoder_0.current_state[2] ),
    .A2(_02435_),
    .ZN(_02456_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _06778_ (.A1(_02435_),
    .A2(_02433_),
    .Z(_02457_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06779_ (.A1(_02456_),
    .A2(_02457_),
    .ZN(_02458_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06780_ (.I(\soc.rom_encoder_0.initializing_step[0] ),
    .Z(_02459_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06781_ (.A1(_02459_),
    .A2(_02449_),
    .ZN(_02460_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06782_ (.A1(_02458_),
    .A2(_02460_),
    .Z(_02461_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _06783_ (.A1(\soc.rom_encoder_0.output_bits_left[4] ),
    .A2(_02440_),
    .Z(_02462_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06784_ (.I(_02462_),
    .Z(_02463_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06785_ (.A1(_02463_),
    .A2(_02458_),
    .ZN(_02464_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06786_ (.A1(\soc.rom_encoder_0.output_buffer[17] ),
    .A2(_02463_),
    .B1(_02464_),
    .B2(\soc.rom_encoder_0.request_data_out[13] ),
    .ZN(_02465_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06787_ (.A1(_02443_),
    .A2(_02465_),
    .ZN(_02466_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _06788_ (.A1(\soc.rom_encoder_0.output_buffer[17] ),
    .A2(_02455_),
    .B(_02461_),
    .C(_02466_),
    .ZN(_02467_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06789_ (.A1(net65),
    .A2(_02453_),
    .ZN(_02468_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _06790_ (.A1(_02453_),
    .A2(_02467_),
    .B(_02468_),
    .C(_01381_),
    .ZN(_00215_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06791_ (.A1(\soc.rom_encoder_0.output_buffer[18] ),
    .A2(_02463_),
    .B1(_02464_),
    .B2(\soc.rom_encoder_0.request_data_out[14] ),
    .ZN(_02469_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06792_ (.A1(_02443_),
    .A2(_02469_),
    .ZN(_02470_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _06793_ (.A1(\soc.rom_encoder_0.output_buffer[18] ),
    .A2(_02455_),
    .B(_02470_),
    .C(_02461_),
    .ZN(_02471_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06794_ (.A1(net66),
    .A2(_02453_),
    .ZN(_02472_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _06795_ (.A1(_02453_),
    .A2(_02471_),
    .B(_02472_),
    .C(_01381_),
    .ZN(_00216_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06796_ (.A1(\soc.rom_encoder_0.output_buffer[19] ),
    .A2(_02463_),
    .B1(_02464_),
    .B2(\soc.rom_encoder_0.request_data_out[15] ),
    .ZN(_02473_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06797_ (.A1(_02443_),
    .A2(_02473_),
    .ZN(_02474_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _06798_ (.A1(\soc.rom_encoder_0.output_buffer[19] ),
    .A2(_02455_),
    .B(_02474_),
    .C(_02461_),
    .ZN(_02475_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06799_ (.A1(net67),
    .A2(_02453_),
    .ZN(_02476_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _06800_ (.A1(_02453_),
    .A2(_02475_),
    .B(_02476_),
    .C(_01381_),
    .ZN(_00217_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06801_ (.I(\soc.ram_encoder_0.output_bits_left[3] ),
    .ZN(_02477_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06802_ (.A1(_02477_),
    .A2(\soc.ram_encoder_0.output_bits_left[2] ),
    .ZN(_02478_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06803_ (.A1(\soc.ram_encoder_0.output_bits_left[4] ),
    .A2(_02478_),
    .ZN(_02479_));
 gf180mcu_fd_sc_mcu7t5v0__inv_3 _06804_ (.I(\soc.ram_encoder_0.current_state[2] ),
    .ZN(_02480_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06805_ (.I(\soc.ram_encoder_0.current_state[1] ),
    .Z(_02481_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06806_ (.I(\soc.ram_encoder_0.current_state[0] ),
    .Z(_02482_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06807_ (.A1(_02480_),
    .A2(_02481_),
    .A3(_02482_),
    .ZN(_02483_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06808_ (.I(\soc.ram_encoder_0.current_state[2] ),
    .Z(_02484_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _06809_ (.I(_02482_),
    .ZN(_02485_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06810_ (.A1(_02481_),
    .A2(_02485_),
    .ZN(_02486_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06811_ (.A1(_02484_),
    .A2(_02486_),
    .ZN(_02487_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06812_ (.A1(\soc.ram_encoder_0.request_write ),
    .A2(_02483_),
    .B(_02487_),
    .ZN(_02488_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06813_ (.A1(_02479_),
    .A2(_02488_),
    .ZN(_02489_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06814_ (.A1(_02481_),
    .A2(_02482_),
    .ZN(_02490_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _06815_ (.I(\soc.ram_encoder_0.current_state[1] ),
    .ZN(_02491_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06816_ (.A1(_02480_),
    .A2(_02491_),
    .ZN(_02492_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06817_ (.A1(_02490_),
    .A2(_02492_),
    .ZN(_02493_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _06818_ (.A1(_01379_),
    .A2(\soc.ram_encoder_0.toggled_sram_sck ),
    .A3(_02489_),
    .A4(_02493_),
    .ZN(_02494_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06819_ (.A1(\soc.ram_encoder_0.output_bits_left[3] ),
    .A2(_02494_),
    .ZN(_02495_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06820_ (.A1(\soc.ram_encoder_0.output_bits_left[3] ),
    .A2(\soc.ram_encoder_0.output_bits_left[2] ),
    .ZN(_02496_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06821_ (.A1(_02484_),
    .A2(_02481_),
    .ZN(_02497_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06822_ (.A1(_02491_),
    .A2(_02485_),
    .ZN(_02498_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06823_ (.A1(_02484_),
    .A2(_02481_),
    .ZN(_02499_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06824_ (.A1(_02498_),
    .A2(_02499_),
    .ZN(_02500_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _06825_ (.A1(\soc.ram_encoder_0.output_bits_left[4] ),
    .A2(_02496_),
    .B(_02497_),
    .C(_02500_),
    .ZN(_02501_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _06826_ (.A1(\soc.ram_encoder_0.output_bits_left[4] ),
    .A2(_02495_),
    .B1(_02501_),
    .B2(_02494_),
    .ZN(_02502_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06827_ (.I(_02502_),
    .ZN(_00218_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _06828_ (.A1(\soc.ram_encoder_0.output_bits_left[4] ),
    .A2(_02478_),
    .Z(_02503_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06829_ (.A1(_02481_),
    .A2(_02485_),
    .ZN(_02504_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _06830_ (.A1(_02484_),
    .A2(_02503_),
    .A3(_02504_),
    .ZN(_02505_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06831_ (.I(_02505_),
    .Z(_02506_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06832_ (.A1(_02477_),
    .A2(\soc.ram_encoder_0.output_bits_left[2] ),
    .Z(_02507_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _06833_ (.A1(_02500_),
    .A2(_02497_),
    .A3(_02506_),
    .A4(_02507_),
    .ZN(_02508_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06834_ (.A1(\soc.ram_encoder_0.output_bits_left[3] ),
    .A2(_02494_),
    .ZN(_02509_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06835_ (.A1(_02494_),
    .A2(_02508_),
    .B(_02509_),
    .ZN(_00219_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06836_ (.A1(_02482_),
    .A2(_02497_),
    .Z(_02510_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _06837_ (.A1(\soc.ram_encoder_0.output_bits_left[2] ),
    .A2(_02494_),
    .A3(_02510_),
    .Z(_02511_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06838_ (.A1(\soc.ram_encoder_0.output_bits_left[2] ),
    .A2(_02494_),
    .ZN(_02512_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06839_ (.A1(_02511_),
    .A2(_02512_),
    .ZN(_00220_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _06840_ (.A1(_01379_),
    .A2(_02456_),
    .A3(_02448_),
    .ZN(_02513_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06841_ (.A1(\soc.rom_encoder_0.output_bits_left[3] ),
    .A2(_02513_),
    .ZN(_02514_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06842_ (.A1(_02434_),
    .A2(_02435_),
    .ZN(_02515_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06843_ (.A1(\soc.rom_encoder_0.output_bits_left[3] ),
    .A2(\soc.rom_encoder_0.output_bits_left[2] ),
    .ZN(_02516_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06844_ (.A1(_02445_),
    .A2(_02515_),
    .B1(_02516_),
    .B2(\soc.rom_encoder_0.output_bits_left[4] ),
    .ZN(_02517_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _06845_ (.A1(\soc.rom_encoder_0.output_bits_left[4] ),
    .A2(_02514_),
    .B1(_02517_),
    .B2(_02513_),
    .ZN(_02518_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06846_ (.I(_02518_),
    .ZN(_00221_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _06847_ (.A1(_02454_),
    .A2(_02515_),
    .A3(_02463_),
    .ZN(_02519_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06848_ (.I(_02519_),
    .Z(_02520_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06849_ (.A1(_02439_),
    .A2(\soc.rom_encoder_0.output_bits_left[2] ),
    .Z(_02521_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _06850_ (.A1(_02445_),
    .A2(_02515_),
    .B(_02520_),
    .C(_02521_),
    .ZN(_02522_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06851_ (.A1(\soc.rom_encoder_0.output_bits_left[3] ),
    .A2(_02513_),
    .ZN(_02523_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06852_ (.A1(_02513_),
    .A2(_02522_),
    .B(_02523_),
    .ZN(_00222_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06853_ (.A1(_02434_),
    .A2(_02454_),
    .ZN(_02524_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06854_ (.A1(_02435_),
    .A2(_02524_),
    .ZN(_02525_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _06855_ (.A1(\soc.rom_encoder_0.output_bits_left[2] ),
    .A2(_02513_),
    .A3(_02525_),
    .Z(_02526_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06856_ (.A1(\soc.rom_encoder_0.output_bits_left[2] ),
    .A2(_02513_),
    .ZN(_02527_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06857_ (.A1(_02526_),
    .A2(_02527_),
    .ZN(_00223_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06858_ (.I(\soc.cpu.AReg.data[15] ),
    .ZN(_02528_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06859_ (.A1(_01822_),
    .A2(_01825_),
    .ZN(_02529_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06860_ (.A1(_01669_),
    .A2(_02529_),
    .ZN(_02530_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _06861_ (.A1(_01831_),
    .A2(_02530_),
    .Z(_02531_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06862_ (.A1(_01618_),
    .A2(\soc.cpu.AReg.data[15] ),
    .B1(_01718_),
    .B2(\soc.ram_data_out[15] ),
    .ZN(_02532_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06863_ (.A1(_01717_),
    .A2(_02532_),
    .ZN(_02533_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06864_ (.A1(_01705_),
    .A2(_02533_),
    .Z(_02534_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06865_ (.A1(_01670_),
    .A2(\soc.cpu.ALU.x[15] ),
    .ZN(_02535_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06866_ (.A1(_01702_),
    .A2(_02535_),
    .Z(_02536_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06867_ (.A1(_01682_),
    .A2(_02534_),
    .B(_02536_),
    .ZN(_02537_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06868_ (.A1(_02534_),
    .A2(_02536_),
    .B(_02537_),
    .ZN(_02538_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _06869_ (.A1(_01654_),
    .A2(_02531_),
    .A3(_02538_),
    .Z(_02539_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _06870_ (.A1(_02528_),
    .A2(_01592_),
    .B1(_02539_),
    .B2(_01555_),
    .ZN(_00224_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06871_ (.A1(_02438_),
    .A2(_02452_),
    .ZN(_02540_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06872_ (.A1(_01379_),
    .A2(_02540_),
    .ZN(_02541_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06873_ (.I(_02541_),
    .Z(_02542_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _06874_ (.A1(_01380_),
    .A2(_02540_),
    .A3(_02519_),
    .Z(_02543_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06875_ (.A1(\soc.rom_encoder_0.output_buffer[4] ),
    .A2(_02542_),
    .B1(_02543_),
    .B2(\soc.rom_encoder_0.request_address[3] ),
    .ZN(_02544_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06876_ (.I(_02544_),
    .ZN(_00225_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06877_ (.A1(\soc.rom_encoder_0.output_buffer[3] ),
    .A2(_02542_),
    .B1(_02543_),
    .B2(\soc.rom_encoder_0.request_address[2] ),
    .ZN(_02545_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06878_ (.I(_02545_),
    .ZN(_00226_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06879_ (.A1(\soc.rom_encoder_0.output_buffer[2] ),
    .A2(_02542_),
    .B1(_02543_),
    .B2(\soc.rom_encoder_0.request_address[1] ),
    .ZN(_02546_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06880_ (.I(_02546_),
    .ZN(_00227_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06881_ (.A1(\soc.rom_encoder_0.output_buffer[1] ),
    .A2(_02542_),
    .B1(_02543_),
    .B2(\soc.rom_encoder_0.request_address[0] ),
    .ZN(_02547_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06882_ (.I(_02547_),
    .ZN(_00228_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06883_ (.A1(_02482_),
    .A2(_02492_),
    .ZN(_02548_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _06884_ (.A1(\soc.ram_encoder_0.initializing_step[4] ),
    .A2(\soc.ram_encoder_0.initializing_step[3] ),
    .Z(_02549_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _06885_ (.A1(\soc.ram_encoder_0.initializing_step[2] ),
    .A2(\soc.ram_encoder_0.initializing_step[1] ),
    .A3(_02549_),
    .ZN(_02550_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06886_ (.A1(_02482_),
    .A2(_02550_),
    .ZN(_02551_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06887_ (.A1(_02492_),
    .A2(_02551_),
    .ZN(_02552_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _06888_ (.A1(\soc.ram_encoder_0.toggled_sram_sck ),
    .A2(_02489_),
    .A3(_02498_),
    .A4(_02552_),
    .ZN(_02553_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _06889_ (.I(_02553_),
    .ZN(_02554_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _06890_ (.A1(_01379_),
    .A2(_02548_),
    .A3(_02554_),
    .ZN(_02555_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06891_ (.I(_02555_),
    .Z(_02556_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06892_ (.A1(\soc.ram_encoder_0.request_address[3] ),
    .A2(_02506_),
    .ZN(_02557_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06893_ (.I(_02555_),
    .Z(_02558_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06894_ (.A1(\soc.ram_encoder_0.output_buffer[4] ),
    .A2(_02558_),
    .ZN(_02559_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06895_ (.A1(_02556_),
    .A2(_02557_),
    .B(_02559_),
    .ZN(_00229_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06896_ (.A1(\soc.ram_encoder_0.request_address[2] ),
    .A2(_02506_),
    .ZN(_02560_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06897_ (.A1(\soc.ram_encoder_0.output_buffer[3] ),
    .A2(_02558_),
    .ZN(_02561_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06898_ (.A1(_02556_),
    .A2(_02560_),
    .B(_02561_),
    .ZN(_00230_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06899_ (.A1(\soc.ram_encoder_0.request_address[1] ),
    .A2(_02506_),
    .ZN(_02562_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06900_ (.I(_02555_),
    .Z(_02563_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06901_ (.A1(\soc.ram_encoder_0.output_buffer[2] ),
    .A2(_02563_),
    .ZN(_02564_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06902_ (.A1(_02556_),
    .A2(_02562_),
    .B(_02564_),
    .ZN(_00231_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06903_ (.A1(\soc.ram_encoder_0.request_address[0] ),
    .A2(_02506_),
    .ZN(_02565_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06904_ (.A1(\soc.ram_encoder_0.output_buffer[1] ),
    .A2(_02563_),
    .ZN(_02566_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06905_ (.A1(_02556_),
    .A2(_02565_),
    .B(_02566_),
    .ZN(_00232_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06906_ (.I(_00004_),
    .Z(_02567_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06907_ (.I(_02567_),
    .Z(_02568_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _06908_ (.I(_00002_),
    .ZN(_02569_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06909_ (.I(_02569_),
    .Z(_02570_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06910_ (.I(_02570_),
    .Z(_02571_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06911_ (.I(_00000_),
    .Z(_02572_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06912_ (.I(_02572_),
    .Z(_02573_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06913_ (.I(_02573_),
    .Z(_02574_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 _06914_ (.I(_02574_),
    .Z(_02575_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06915_ (.I(_00001_),
    .Z(_02576_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06916_ (.I(_02576_),
    .Z(_02577_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06917_ (.I(_02577_),
    .Z(_02578_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06918_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[12][0] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[13][0] ),
    .I2(\soc.spi_video_ram_1.write_fifo.fifo_mem[14][0] ),
    .I3(\soc.spi_video_ram_1.write_fifo.fifo_mem[15][0] ),
    .S0(_02575_),
    .S1(_02578_),
    .Z(_02579_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06919_ (.A1(_02571_),
    .A2(_02579_),
    .ZN(_02580_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06920_ (.I(_00002_),
    .Z(_02581_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06921_ (.I(_02581_),
    .Z(_02582_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06922_ (.I(_02582_),
    .Z(_02583_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06923_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[8][0] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[9][0] ),
    .I2(\soc.spi_video_ram_1.write_fifo.fifo_mem[10][0] ),
    .I3(\soc.spi_video_ram_1.write_fifo.fifo_mem[11][0] ),
    .S0(_02575_),
    .S1(_02578_),
    .Z(_02584_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06924_ (.I(_00003_),
    .Z(_02585_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06925_ (.I(_02585_),
    .Z(_02586_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06926_ (.A1(_02583_),
    .A2(_02584_),
    .B(_02586_),
    .ZN(_02587_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06927_ (.I(_02581_),
    .Z(_02588_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06928_ (.I(_02588_),
    .Z(_02589_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06929_ (.I(_02572_),
    .Z(_02590_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06930_ (.I(_02590_),
    .Z(_02591_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06931_ (.I(_02576_),
    .Z(_02592_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06932_ (.I(_02592_),
    .Z(_02593_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06933_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[0][0] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[1][0] ),
    .I2(\soc.spi_video_ram_1.write_fifo.fifo_mem[2][0] ),
    .I3(\soc.spi_video_ram_1.write_fifo.fifo_mem[3][0] ),
    .S0(_02591_),
    .S1(_02593_),
    .Z(_02594_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06934_ (.A1(_02589_),
    .A2(_02594_),
    .ZN(_02595_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06935_ (.I(_02570_),
    .Z(_02596_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06936_ (.I(_02590_),
    .Z(_02597_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06937_ (.I(_02592_),
    .Z(_02598_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06938_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[4][0] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[5][0] ),
    .I2(\soc.spi_video_ram_1.write_fifo.fifo_mem[6][0] ),
    .I3(\soc.spi_video_ram_1.write_fifo.fifo_mem[7][0] ),
    .S0(_02597_),
    .S1(_02598_),
    .Z(_02599_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06939_ (.I(_00003_),
    .ZN(_02600_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06940_ (.I(_02600_),
    .Z(_02601_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06941_ (.I(_02601_),
    .Z(_02602_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06942_ (.A1(_02596_),
    .A2(_02599_),
    .B(_02602_),
    .ZN(_02603_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _06943_ (.A1(_02580_),
    .A2(_02587_),
    .B1(_02595_),
    .B2(_02603_),
    .ZN(_02604_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06944_ (.A1(_02568_),
    .A2(_02604_),
    .ZN(_02605_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06945_ (.I(_01391_),
    .Z(_02606_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06946_ (.I(_02590_),
    .Z(_02607_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06947_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[28][0] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[29][0] ),
    .I2(\soc.spi_video_ram_1.write_fifo.fifo_mem[30][0] ),
    .I3(\soc.spi_video_ram_1.write_fifo.fifo_mem[31][0] ),
    .S0(_02607_),
    .S1(_02578_),
    .Z(_02608_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06948_ (.A1(_02596_),
    .A2(_02608_),
    .ZN(_02609_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06949_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[24][0] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[25][0] ),
    .I2(\soc.spi_video_ram_1.write_fifo.fifo_mem[26][0] ),
    .I3(\soc.spi_video_ram_1.write_fifo.fifo_mem[27][0] ),
    .S0(_02607_),
    .S1(_02578_),
    .Z(_02610_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06950_ (.A1(_02583_),
    .A2(_02610_),
    .B(_02586_),
    .ZN(_02611_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06951_ (.I(_02572_),
    .Z(_02612_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 _06952_ (.I(_02612_),
    .Z(_02613_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06953_ (.I(_02592_),
    .Z(_02614_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06954_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[16][0] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[17][0] ),
    .I2(\soc.spi_video_ram_1.write_fifo.fifo_mem[18][0] ),
    .I3(\soc.spi_video_ram_1.write_fifo.fifo_mem[19][0] ),
    .S0(_02613_),
    .S1(_02614_),
    .Z(_02615_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06955_ (.A1(_02589_),
    .A2(_02615_),
    .ZN(_02616_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06956_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[20][0] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[21][0] ),
    .I2(\soc.spi_video_ram_1.write_fifo.fifo_mem[22][0] ),
    .I3(\soc.spi_video_ram_1.write_fifo.fifo_mem[23][0] ),
    .S0(_02591_),
    .S1(_02593_),
    .Z(_02617_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06957_ (.I(_02601_),
    .Z(_02618_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06958_ (.A1(_02596_),
    .A2(_02617_),
    .B(_02618_),
    .ZN(_02619_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06959_ (.I(_00004_),
    .Z(_02620_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _06960_ (.A1(_02609_),
    .A2(_02611_),
    .B1(_02616_),
    .B2(_02619_),
    .C(_02620_),
    .ZN(_02621_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06961_ (.A1(_02606_),
    .A2(_02621_),
    .ZN(_02622_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06962_ (.A1(_02054_),
    .A2(_02057_),
    .ZN(_02623_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _06963_ (.A1(\soc.spi_video_ram_1.state_sram_clk_counter[1] ),
    .A2(_01391_),
    .Z(_02624_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06964_ (.A1(_01419_),
    .A2(_02624_),
    .ZN(_02625_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _06965_ (.A1(_02623_),
    .A2(_02625_),
    .Z(_02626_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06966_ (.A1(_01411_),
    .A2(_02626_),
    .Z(_02627_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06967_ (.A1(_02605_),
    .A2(_02622_),
    .B(_02627_),
    .ZN(_02628_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _06968_ (.I(_02624_),
    .ZN(_02629_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06969_ (.A1(_01428_),
    .A2(\soc.spi_video_ram_1.current_state[0] ),
    .ZN(_02630_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _06970_ (.A1(\soc.spi_video_ram_1.current_state[4] ),
    .A2(_01417_),
    .B(_01391_),
    .ZN(_02631_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_4 _06971_ (.A1(\soc.spi_video_ram_1.current_state[0] ),
    .A2(_01411_),
    .B1(_02629_),
    .B2(_02630_),
    .C(_02631_),
    .ZN(_02632_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _06972_ (.A1(_01378_),
    .A2(_02632_),
    .ZN(_02633_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06973_ (.I0(\soc.spi_video_ram_1.output_buffer[23] ),
    .I1(_02628_),
    .S(_02633_),
    .Z(_02634_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06974_ (.I(_02634_),
    .Z(_00233_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06975_ (.I(_02612_),
    .Z(_02635_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06976_ (.I(_02592_),
    .Z(_02636_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06977_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[8][1] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[9][1] ),
    .I2(\soc.spi_video_ram_1.write_fifo.fifo_mem[10][1] ),
    .I3(\soc.spi_video_ram_1.write_fifo.fifo_mem[11][1] ),
    .S0(_02635_),
    .S1(_02636_),
    .Z(_02637_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06978_ (.A1(_02583_),
    .A2(_02637_),
    .ZN(_02638_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06979_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[12][1] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[13][1] ),
    .I2(\soc.spi_video_ram_1.write_fifo.fifo_mem[14][1] ),
    .I3(\soc.spi_video_ram_1.write_fifo.fifo_mem[15][1] ),
    .S0(_02607_),
    .S1(_02636_),
    .Z(_02639_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06980_ (.I(_02585_),
    .Z(_02640_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06981_ (.A1(_02571_),
    .A2(_02639_),
    .B(_02640_),
    .ZN(_02641_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06982_ (.I(_00002_),
    .Z(_02642_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06983_ (.I(_02642_),
    .Z(_02643_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06984_ (.I(_02572_),
    .Z(_02644_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06985_ (.I(_02644_),
    .Z(_02645_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06986_ (.I(_02576_),
    .Z(_02646_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06987_ (.I(_02646_),
    .Z(_02647_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06988_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[0][1] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[1][1] ),
    .I2(\soc.spi_video_ram_1.write_fifo.fifo_mem[2][1] ),
    .I3(\soc.spi_video_ram_1.write_fifo.fifo_mem[3][1] ),
    .S0(_02645_),
    .S1(_02647_),
    .Z(_02648_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06989_ (.A1(_02643_),
    .A2(_02648_),
    .ZN(_02649_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06990_ (.I(_02569_),
    .Z(_02650_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06991_ (.I(_02612_),
    .Z(_02651_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06992_ (.I(_02592_),
    .Z(_02652_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06993_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[4][1] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[5][1] ),
    .I2(\soc.spi_video_ram_1.write_fifo.fifo_mem[6][1] ),
    .I3(\soc.spi_video_ram_1.write_fifo.fifo_mem[7][1] ),
    .S0(_02651_),
    .S1(_02652_),
    .Z(_02653_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06994_ (.A1(_02650_),
    .A2(_02653_),
    .B(_02618_),
    .ZN(_02654_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _06995_ (.I(_00004_),
    .ZN(_02655_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06996_ (.I(_02655_),
    .Z(_02656_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _06997_ (.A1(_02638_),
    .A2(_02641_),
    .B1(_02649_),
    .B2(_02654_),
    .C(_02656_),
    .ZN(_02657_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _06998_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[28][1] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[29][1] ),
    .I2(\soc.spi_video_ram_1.write_fifo.fifo_mem[30][1] ),
    .I3(\soc.spi_video_ram_1.write_fifo.fifo_mem[31][1] ),
    .S0(_02635_),
    .S1(_02636_),
    .Z(_02658_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06999_ (.A1(_02596_),
    .A2(_02658_),
    .ZN(_02659_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _07000_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[24][1] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[25][1] ),
    .I2(\soc.spi_video_ram_1.write_fifo.fifo_mem[26][1] ),
    .I3(\soc.spi_video_ram_1.write_fifo.fifo_mem[27][1] ),
    .S0(_02635_),
    .S1(_02636_),
    .Z(_02660_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07001_ (.A1(_02583_),
    .A2(_02660_),
    .B(_02640_),
    .ZN(_02661_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _07002_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[16][1] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[17][1] ),
    .I2(\soc.spi_video_ram_1.write_fifo.fifo_mem[18][1] ),
    .I3(\soc.spi_video_ram_1.write_fifo.fifo_mem[19][1] ),
    .S0(_02645_),
    .S1(_02614_),
    .Z(_02662_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07003_ (.A1(_02589_),
    .A2(_02662_),
    .ZN(_02663_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _07004_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[20][1] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[21][1] ),
    .I2(\soc.spi_video_ram_1.write_fifo.fifo_mem[22][1] ),
    .I3(\soc.spi_video_ram_1.write_fifo.fifo_mem[23][1] ),
    .S0(_02651_),
    .S1(_02593_),
    .Z(_02664_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07005_ (.A1(_02650_),
    .A2(_02664_),
    .B(_02618_),
    .ZN(_02665_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _07006_ (.A1(_02659_),
    .A2(_02661_),
    .B1(_02663_),
    .B2(_02665_),
    .C(_02620_),
    .ZN(_02666_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07007_ (.A1(_02606_),
    .A2(_02657_),
    .A3(_02666_),
    .ZN(_02667_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07008_ (.A1(_02627_),
    .A2(_02667_),
    .ZN(_02668_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07009_ (.I0(\soc.spi_video_ram_1.output_buffer[22] ),
    .I1(_02668_),
    .S(_02633_),
    .Z(_02669_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07010_ (.I(_02669_),
    .Z(_00234_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07011_ (.I(\soc.spi_video_ram_1.output_buffer[21] ),
    .ZN(_02670_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07012_ (.A1(_02630_),
    .A2(_02631_),
    .ZN(_02671_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07013_ (.A1(_02624_),
    .A2(_02671_),
    .ZN(_02672_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07014_ (.A1(\soc.spi_video_ram_1.current_state[0] ),
    .A2(_01411_),
    .ZN(_02673_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07015_ (.A1(net18),
    .A2(_02673_),
    .ZN(_02674_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07016_ (.A1(_02672_),
    .A2(_02674_),
    .ZN(_02675_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07017_ (.I(_02675_),
    .Z(_02676_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07018_ (.I(\soc.spi_video_ram_1.current_state[1] ),
    .Z(_02677_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07019_ (.I(_02643_),
    .Z(_02678_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _07020_ (.I(_02572_),
    .Z(_02679_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _07021_ (.I(_02679_),
    .Z(_02680_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _07022_ (.I(_02680_),
    .Z(_02681_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _07023_ (.I(_02598_),
    .Z(_02682_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _07024_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[8][2] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[9][2] ),
    .I2(\soc.spi_video_ram_1.write_fifo.fifo_mem[10][2] ),
    .I3(\soc.spi_video_ram_1.write_fifo.fifo_mem[11][2] ),
    .S0(_02681_),
    .S1(_02682_),
    .Z(_02683_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07025_ (.A1(_02678_),
    .A2(_02683_),
    .ZN(_02684_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07026_ (.I(_02596_),
    .Z(_02685_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _07027_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[12][2] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[13][2] ),
    .I2(\soc.spi_video_ram_1.write_fifo.fifo_mem[14][2] ),
    .I3(\soc.spi_video_ram_1.write_fifo.fifo_mem[15][2] ),
    .S0(_02681_),
    .S1(_02682_),
    .Z(_02686_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07028_ (.A1(_02685_),
    .A2(_02686_),
    .B(_02586_),
    .ZN(_02687_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _07029_ (.I(_02644_),
    .Z(_02688_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _07030_ (.I(_02688_),
    .Z(_02689_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07031_ (.I(_02576_),
    .Z(_02690_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07032_ (.I(_02690_),
    .Z(_02691_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _07033_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[0][2] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[1][2] ),
    .I2(\soc.spi_video_ram_1.write_fifo.fifo_mem[2][2] ),
    .I3(\soc.spi_video_ram_1.write_fifo.fifo_mem[3][2] ),
    .S0(_02689_),
    .S1(_02691_),
    .Z(_02692_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07034_ (.I(_02598_),
    .Z(_02693_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07035_ (.I(_02572_),
    .ZN(_02694_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07036_ (.I(_02694_),
    .Z(_02695_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07037_ (.I(_02695_),
    .Z(_02696_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07038_ (.I(_02696_),
    .Z(_02697_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _07039_ (.A1(_02597_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[4][2] ),
    .Z(_02698_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07040_ (.A1(_02697_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[5][2] ),
    .B(_02698_),
    .ZN(_02699_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 _07041_ (.I(_02644_),
    .Z(_02700_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _07042_ (.I(_02700_),
    .Z(_02701_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07043_ (.A1(_02701_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[6][2] ),
    .ZN(_02702_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07044_ (.I(_02694_),
    .Z(_02703_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07045_ (.I(_02703_),
    .Z(_02704_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07046_ (.A1(_02704_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[7][2] ),
    .B(_02691_),
    .ZN(_02705_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07047_ (.I(_00002_),
    .Z(_02706_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07048_ (.I(_02706_),
    .Z(_02707_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _07049_ (.A1(_02693_),
    .A2(_02699_),
    .B1(_02702_),
    .B2(_02705_),
    .C(_02707_),
    .ZN(_02708_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07050_ (.A1(_02583_),
    .A2(_02692_),
    .B(_02708_),
    .C(_02602_),
    .ZN(_02709_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07051_ (.I(_02655_),
    .Z(_02710_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07052_ (.A1(_02684_),
    .A2(_02687_),
    .B(_02709_),
    .C(_02710_),
    .ZN(_02711_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _07053_ (.I(_02644_),
    .Z(_02712_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _07054_ (.I(_02712_),
    .Z(_02713_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _07055_ (.I(_02598_),
    .Z(_02714_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _07056_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[16][2] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[17][2] ),
    .I2(\soc.spi_video_ram_1.write_fifo.fifo_mem[18][2] ),
    .I3(\soc.spi_video_ram_1.write_fifo.fifo_mem[19][2] ),
    .S0(_02713_),
    .S1(_02714_),
    .Z(_02715_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07057_ (.A1(_02678_),
    .A2(_02715_),
    .ZN(_02716_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _07058_ (.I(_02712_),
    .Z(_02717_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _07059_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[20][2] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[21][2] ),
    .I2(\soc.spi_video_ram_1.write_fifo.fifo_mem[22][2] ),
    .I3(\soc.spi_video_ram_1.write_fifo.fifo_mem[23][2] ),
    .S0(_02717_),
    .S1(_02714_),
    .Z(_02718_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07060_ (.I(_02601_),
    .Z(_02719_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07061_ (.I(_02719_),
    .Z(_02720_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07062_ (.A1(_02685_),
    .A2(_02718_),
    .B(_02720_),
    .ZN(_02721_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07063_ (.I(_02646_),
    .Z(_02722_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07064_ (.I(_02722_),
    .Z(_02723_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _07065_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[24][2] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[25][2] ),
    .I2(\soc.spi_video_ram_1.write_fifo.fifo_mem[26][2] ),
    .I3(\soc.spi_video_ram_1.write_fifo.fifo_mem[27][2] ),
    .S0(_02689_),
    .S1(_02723_),
    .Z(_02724_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07066_ (.A1(_02697_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[31][2] ),
    .ZN(_02725_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 _07067_ (.I(_02607_),
    .Z(_02726_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07068_ (.A1(_02726_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[30][2] ),
    .B(_02691_),
    .ZN(_02727_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _07069_ (.A1(_02651_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[29][2] ),
    .Z(_02728_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07070_ (.A1(_02704_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[28][2] ),
    .B(_02728_),
    .ZN(_02729_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _07071_ (.A1(_02725_),
    .A2(_02727_),
    .B1(_02729_),
    .B2(_02693_),
    .C(_02707_),
    .ZN(_02730_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07072_ (.A1(_02583_),
    .A2(_02724_),
    .B(_02730_),
    .C(_02586_),
    .ZN(_02731_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07073_ (.A1(_02716_),
    .A2(_02721_),
    .B(_02731_),
    .C(_02568_),
    .ZN(_02732_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _07074_ (.A1(_02677_),
    .A2(_02606_),
    .A3(_02711_),
    .A4(_02732_),
    .ZN(_02733_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07075_ (.I(_02674_),
    .ZN(_00830_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _07076_ (.A1(_02624_),
    .A2(_02671_),
    .B(_00830_),
    .ZN(_02734_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _07077_ (.A1(_01409_),
    .A2(_01411_),
    .A3(_02734_),
    .A4(_02626_),
    .Z(_02735_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07078_ (.A1(_02670_),
    .A2(_02676_),
    .B1(_02733_),
    .B2(_02735_),
    .ZN(_00235_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07079_ (.I(_02643_),
    .Z(_02736_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _07080_ (.I(_02636_),
    .Z(_02737_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _07081_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[0][3] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[1][3] ),
    .I2(\soc.spi_video_ram_1.write_fifo.fifo_mem[2][3] ),
    .I3(\soc.spi_video_ram_1.write_fifo.fifo_mem[3][3] ),
    .S0(_02713_),
    .S1(_02737_),
    .Z(_02738_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07082_ (.A1(_02726_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[4][3] ),
    .ZN(_02739_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _07083_ (.I(_02576_),
    .ZN(_02740_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07084_ (.I(_02740_),
    .Z(_02741_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07085_ (.I(_02741_),
    .Z(_02742_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07086_ (.A1(_02697_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[5][3] ),
    .B(_02742_),
    .ZN(_02743_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07087_ (.I(_02590_),
    .Z(_02744_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _07088_ (.A1(_02744_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[6][3] ),
    .Z(_02745_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07089_ (.A1(_02697_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[7][3] ),
    .B(_02745_),
    .C(_02723_),
    .ZN(_02746_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07090_ (.A1(_02739_),
    .A2(_02743_),
    .B(_02589_),
    .C(_02746_),
    .ZN(_02747_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07091_ (.A1(_02736_),
    .A2(_02738_),
    .B(_02747_),
    .C(_02720_),
    .ZN(_02748_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _07092_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[8][3] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[9][3] ),
    .I2(\soc.spi_video_ram_1.write_fifo.fifo_mem[10][3] ),
    .I3(\soc.spi_video_ram_1.write_fifo.fifo_mem[11][3] ),
    .S0(_02713_),
    .S1(_02714_),
    .Z(_02749_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07093_ (.A1(_02697_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[15][3] ),
    .ZN(_02750_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07094_ (.A1(_02726_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[14][3] ),
    .B(_02714_),
    .ZN(_02751_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07095_ (.I(_02574_),
    .Z(_02752_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _07096_ (.A1(_02752_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[13][3] ),
    .Z(_02753_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07097_ (.A1(_02697_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[12][3] ),
    .B(_02753_),
    .ZN(_02754_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _07098_ (.A1(_02750_),
    .A2(_02751_),
    .B1(_02754_),
    .B2(_02693_),
    .C(_02643_),
    .ZN(_02755_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07099_ (.A1(_02678_),
    .A2(_02749_),
    .B(_02755_),
    .C(_02586_),
    .ZN(_02756_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07100_ (.A1(_02710_),
    .A2(_02748_),
    .A3(_02756_),
    .ZN(_02757_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _07101_ (.I(_02598_),
    .Z(_02758_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _07102_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[16][3] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[17][3] ),
    .I2(\soc.spi_video_ram_1.write_fifo.fifo_mem[18][3] ),
    .I3(\soc.spi_video_ram_1.write_fifo.fifo_mem[19][3] ),
    .S0(_02681_),
    .S1(_02758_),
    .Z(_02759_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07103_ (.A1(_02678_),
    .A2(_02759_),
    .ZN(_02760_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _07104_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[20][3] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[21][3] ),
    .I2(\soc.spi_video_ram_1.write_fifo.fifo_mem[22][3] ),
    .I3(\soc.spi_video_ram_1.write_fifo.fifo_mem[23][3] ),
    .S0(_02717_),
    .S1(_02682_),
    .Z(_02761_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07105_ (.A1(_02685_),
    .A2(_02761_),
    .B(_02720_),
    .ZN(_02762_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 _07106_ (.I(_02644_),
    .Z(_02763_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 _07107_ (.I(_02763_),
    .Z(_02764_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _07108_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[28][3] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[29][3] ),
    .I2(\soc.spi_video_ram_1.write_fifo.fifo_mem[30][3] ),
    .I3(\soc.spi_video_ram_1.write_fifo.fifo_mem[31][3] ),
    .S0(_02764_),
    .S1(_02723_),
    .Z(_02765_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07109_ (.A1(_02571_),
    .A2(_02765_),
    .B(_02586_),
    .ZN(_02766_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07110_ (.I(_02706_),
    .Z(_02767_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07111_ (.I(_02767_),
    .Z(_02768_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _07112_ (.I(_02763_),
    .Z(_02769_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _07113_ (.I(_02652_),
    .Z(_02770_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _07114_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[24][3] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[25][3] ),
    .I2(\soc.spi_video_ram_1.write_fifo.fifo_mem[26][3] ),
    .I3(\soc.spi_video_ram_1.write_fifo.fifo_mem[27][3] ),
    .S0(_02769_),
    .S1(_02770_),
    .Z(_02771_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07115_ (.A1(_02768_),
    .A2(_02771_),
    .ZN(_02772_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _07116_ (.A1(_02760_),
    .A2(_02762_),
    .B1(_02766_),
    .B2(_02772_),
    .C(_02568_),
    .ZN(_02773_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _07117_ (.A1(_02677_),
    .A2(_02606_),
    .A3(_02757_),
    .A4(_02773_),
    .ZN(_02774_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07118_ (.A1(_01534_),
    .A2(_02676_),
    .B1(_02735_),
    .B2(_02774_),
    .ZN(_00236_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _07119_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[0][4] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[1][4] ),
    .I2(\soc.spi_video_ram_1.write_fifo.fifo_mem[2][4] ),
    .I3(\soc.spi_video_ram_1.write_fifo.fifo_mem[3][4] ),
    .S0(_02713_),
    .S1(_02714_),
    .Z(_02775_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07120_ (.A1(_02726_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[4][4] ),
    .ZN(_02776_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07121_ (.A1(_02697_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[5][4] ),
    .B(_02742_),
    .ZN(_02777_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _07122_ (.A1(_02744_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[6][4] ),
    .Z(_02778_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07123_ (.A1(_02697_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[7][4] ),
    .B(_02778_),
    .C(_02723_),
    .ZN(_02779_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07124_ (.A1(_02776_),
    .A2(_02777_),
    .B(_02589_),
    .C(_02779_),
    .ZN(_02780_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07125_ (.A1(_02736_),
    .A2(_02775_),
    .B(_02780_),
    .C(_02602_),
    .ZN(_02781_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _07126_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[8][4] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[9][4] ),
    .I2(\soc.spi_video_ram_1.write_fifo.fifo_mem[10][4] ),
    .I3(\soc.spi_video_ram_1.write_fifo.fifo_mem[11][4] ),
    .S0(_02713_),
    .S1(_02714_),
    .Z(_02782_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _07127_ (.I(_02573_),
    .Z(_02783_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07128_ (.I(_02783_),
    .Z(_02784_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _07129_ (.A1(_02784_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[13][4] ),
    .Z(_02785_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07130_ (.A1(_02697_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[12][4] ),
    .B(_02785_),
    .ZN(_02786_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07131_ (.A1(_02697_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[15][4] ),
    .ZN(_02787_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07132_ (.A1(_02726_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[14][4] ),
    .B(_02770_),
    .ZN(_02788_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _07133_ (.A1(_02693_),
    .A2(_02786_),
    .B1(_02787_),
    .B2(_02788_),
    .C(_02643_),
    .ZN(_02789_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07134_ (.A1(_02678_),
    .A2(_02782_),
    .B(_02789_),
    .C(_02586_),
    .ZN(_02790_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07135_ (.A1(_02710_),
    .A2(_02781_),
    .A3(_02790_),
    .ZN(_02791_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _07136_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[16][4] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[17][4] ),
    .I2(\soc.spi_video_ram_1.write_fifo.fifo_mem[18][4] ),
    .I3(\soc.spi_video_ram_1.write_fifo.fifo_mem[19][4] ),
    .S0(_02681_),
    .S1(_02758_),
    .Z(_02792_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07137_ (.A1(_02678_),
    .A2(_02792_),
    .ZN(_02793_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _07138_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[20][4] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[21][4] ),
    .I2(\soc.spi_video_ram_1.write_fifo.fifo_mem[22][4] ),
    .I3(\soc.spi_video_ram_1.write_fifo.fifo_mem[23][4] ),
    .S0(_02717_),
    .S1(_02682_),
    .Z(_02794_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07139_ (.A1(_02685_),
    .A2(_02794_),
    .B(_02720_),
    .ZN(_02795_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _07140_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[28][4] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[29][4] ),
    .I2(\soc.spi_video_ram_1.write_fifo.fifo_mem[30][4] ),
    .I3(\soc.spi_video_ram_1.write_fifo.fifo_mem[31][4] ),
    .S0(_02689_),
    .S1(_02723_),
    .Z(_02796_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07141_ (.A1(_02571_),
    .A2(_02796_),
    .B(_02586_),
    .ZN(_02797_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _07142_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[24][4] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[25][4] ),
    .I2(\soc.spi_video_ram_1.write_fifo.fifo_mem[26][4] ),
    .I3(\soc.spi_video_ram_1.write_fifo.fifo_mem[27][4] ),
    .S0(_02769_),
    .S1(_02770_),
    .Z(_02798_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07143_ (.A1(_02768_),
    .A2(_02798_),
    .ZN(_02799_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _07144_ (.A1(_02793_),
    .A2(_02795_),
    .B1(_02797_),
    .B2(_02799_),
    .C(_02568_),
    .ZN(_02800_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _07145_ (.A1(_02677_),
    .A2(_02606_),
    .A3(_02791_),
    .A4(_02800_),
    .ZN(_02801_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07146_ (.A1(_01508_),
    .A2(_02676_),
    .B1(_02735_),
    .B2(_02801_),
    .ZN(_00237_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _07147_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[8][5] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[9][5] ),
    .I2(\soc.spi_video_ram_1.write_fifo.fifo_mem[10][5] ),
    .I3(\soc.spi_video_ram_1.write_fifo.fifo_mem[11][5] ),
    .S0(_02635_),
    .S1(_02636_),
    .Z(_02802_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07148_ (.A1(_02583_),
    .A2(_02802_),
    .ZN(_02803_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _07149_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[12][5] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[13][5] ),
    .I2(\soc.spi_video_ram_1.write_fifo.fifo_mem[14][5] ),
    .I3(\soc.spi_video_ram_1.write_fifo.fifo_mem[15][5] ),
    .S0(_02635_),
    .S1(_02636_),
    .Z(_02804_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07150_ (.A1(_02596_),
    .A2(_02804_),
    .B(_02640_),
    .ZN(_02805_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _07151_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[0][5] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[1][5] ),
    .I2(\soc.spi_video_ram_1.write_fifo.fifo_mem[2][5] ),
    .I3(\soc.spi_video_ram_1.write_fifo.fifo_mem[3][5] ),
    .S0(_02700_),
    .S1(_02647_),
    .Z(_02806_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07152_ (.A1(_02643_),
    .A2(_02806_),
    .ZN(_02807_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _07153_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[4][5] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[5][5] ),
    .I2(\soc.spi_video_ram_1.write_fifo.fifo_mem[6][5] ),
    .I3(\soc.spi_video_ram_1.write_fifo.fifo_mem[7][5] ),
    .S0(_02651_),
    .S1(_02652_),
    .Z(_02808_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07154_ (.A1(_02650_),
    .A2(_02808_),
    .B(_02618_),
    .ZN(_02809_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _07155_ (.A1(_02803_),
    .A2(_02805_),
    .B1(_02807_),
    .B2(_02809_),
    .C(_02656_),
    .ZN(_02810_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _07156_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[28][5] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[29][5] ),
    .I2(\soc.spi_video_ram_1.write_fifo.fifo_mem[30][5] ),
    .I3(\soc.spi_video_ram_1.write_fifo.fifo_mem[31][5] ),
    .S0(_02635_),
    .S1(_02636_),
    .Z(_02811_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07157_ (.A1(_02596_),
    .A2(_02811_),
    .ZN(_02812_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _07158_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[24][5] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[25][5] ),
    .I2(\soc.spi_video_ram_1.write_fifo.fifo_mem[26][5] ),
    .I3(\soc.spi_video_ram_1.write_fifo.fifo_mem[27][5] ),
    .S0(_02635_),
    .S1(_02636_),
    .Z(_02813_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07159_ (.A1(_02583_),
    .A2(_02813_),
    .B(_02640_),
    .ZN(_02814_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _07160_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[16][5] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[17][5] ),
    .I2(\soc.spi_video_ram_1.write_fifo.fifo_mem[18][5] ),
    .I3(\soc.spi_video_ram_1.write_fifo.fifo_mem[19][5] ),
    .S0(_02645_),
    .S1(_02647_),
    .Z(_02815_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07161_ (.A1(_02643_),
    .A2(_02815_),
    .ZN(_02816_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _07162_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[20][5] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[21][5] ),
    .I2(\soc.spi_video_ram_1.write_fifo.fifo_mem[22][5] ),
    .I3(\soc.spi_video_ram_1.write_fifo.fifo_mem[23][5] ),
    .S0(_02651_),
    .S1(_02652_),
    .Z(_02817_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07163_ (.A1(_02650_),
    .A2(_02817_),
    .B(_02618_),
    .ZN(_02818_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _07164_ (.A1(_02812_),
    .A2(_02814_),
    .B1(_02816_),
    .B2(_02818_),
    .C(_02620_),
    .ZN(_02819_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07165_ (.A1(_02606_),
    .A2(_02810_),
    .A3(_02819_),
    .ZN(_02820_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07166_ (.A1(_02627_),
    .A2(_02820_),
    .ZN(_02821_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07167_ (.I0(\soc.spi_video_ram_1.output_buffer[18] ),
    .I1(_02821_),
    .S(_02633_),
    .Z(_02822_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07168_ (.I(_02822_),
    .Z(_00238_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _07169_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[16][6] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[17][6] ),
    .I2(\soc.spi_video_ram_1.write_fifo.fifo_mem[18][6] ),
    .I3(\soc.spi_video_ram_1.write_fifo.fifo_mem[19][6] ),
    .S0(_02645_),
    .S1(_02614_),
    .Z(_02823_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07170_ (.A1(_02589_),
    .A2(_02823_),
    .ZN(_02824_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _07171_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[20][6] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[21][6] ),
    .I2(\soc.spi_video_ram_1.write_fifo.fifo_mem[22][6] ),
    .I3(\soc.spi_video_ram_1.write_fifo.fifo_mem[23][6] ),
    .S0(_02645_),
    .S1(_02614_),
    .Z(_02825_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07172_ (.A1(_02650_),
    .A2(_02825_),
    .B(_02719_),
    .ZN(_02826_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _07173_ (.I(_02646_),
    .Z(_02827_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _07174_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[24][6] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[25][6] ),
    .I2(\soc.spi_video_ram_1.write_fifo.fifo_mem[26][6] ),
    .I3(\soc.spi_video_ram_1.write_fifo.fifo_mem[27][6] ),
    .S0(_02763_),
    .S1(_02827_),
    .Z(_02828_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07175_ (.A1(_02767_),
    .A2(_02828_),
    .ZN(_02829_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _07176_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[28][6] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[29][6] ),
    .I2(\soc.spi_video_ram_1.write_fifo.fifo_mem[30][6] ),
    .I3(\soc.spi_video_ram_1.write_fifo.fifo_mem[31][6] ),
    .S0(_02680_),
    .S1(_02722_),
    .Z(_02830_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07177_ (.I(_02585_),
    .Z(_02831_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07178_ (.A1(_02650_),
    .A2(_02830_),
    .B(_02831_),
    .ZN(_02832_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _07179_ (.A1(_02824_),
    .A2(_02826_),
    .B1(_02829_),
    .B2(_02832_),
    .C(_02567_),
    .ZN(_02833_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _07180_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[0][6] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[1][6] ),
    .I2(\soc.spi_video_ram_1.write_fifo.fifo_mem[2][6] ),
    .I3(\soc.spi_video_ram_1.write_fifo.fifo_mem[3][6] ),
    .S0(_02613_),
    .S1(_02652_),
    .Z(_02834_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07181_ (.A1(_02589_),
    .A2(_02834_),
    .ZN(_02835_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _07182_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[4][6] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[5][6] ),
    .I2(\soc.spi_video_ram_1.write_fifo.fifo_mem[6][6] ),
    .I3(\soc.spi_video_ram_1.write_fifo.fifo_mem[7][6] ),
    .S0(_02613_),
    .S1(_02652_),
    .Z(_02836_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07183_ (.A1(_02650_),
    .A2(_02836_),
    .B(_02618_),
    .ZN(_02837_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _07184_ (.I(_02646_),
    .Z(_02838_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _07185_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[12][6] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[13][6] ),
    .I2(\soc.spi_video_ram_1.write_fifo.fifo_mem[14][6] ),
    .I3(\soc.spi_video_ram_1.write_fifo.fifo_mem[15][6] ),
    .S0(_02680_),
    .S1(_02838_),
    .Z(_02839_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07186_ (.A1(_02570_),
    .A2(_02839_),
    .ZN(_02840_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _07187_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[8][6] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[9][6] ),
    .I2(\soc.spi_video_ram_1.write_fifo.fifo_mem[10][6] ),
    .I3(\soc.spi_video_ram_1.write_fifo.fifo_mem[11][6] ),
    .S0(_02680_),
    .S1(_02722_),
    .Z(_02841_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07188_ (.A1(_02643_),
    .A2(_02841_),
    .B(_02831_),
    .ZN(_02842_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _07189_ (.A1(_02835_),
    .A2(_02837_),
    .B1(_02840_),
    .B2(_02842_),
    .C(_02656_),
    .ZN(_02843_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _07190_ (.A1(_02606_),
    .A2(_02833_),
    .A3(_02843_),
    .Z(_02844_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07191_ (.A1(_02629_),
    .A2(_02844_),
    .B(_02677_),
    .ZN(_02845_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07192_ (.A1(_02623_),
    .A2(_02624_),
    .ZN(_02846_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07193_ (.A1(_01419_),
    .A2(_02846_),
    .ZN(_02847_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _07194_ (.A1(_01411_),
    .A2(_02633_),
    .A3(_02847_),
    .Z(_02848_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07195_ (.A1(_01507_),
    .A2(_02676_),
    .B1(_02845_),
    .B2(_02848_),
    .ZN(_00239_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _07196_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[28][7] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[29][7] ),
    .I2(\soc.spi_video_ram_1.write_fifo.fifo_mem[30][7] ),
    .I3(\soc.spi_video_ram_1.write_fifo.fifo_mem[31][7] ),
    .S0(_02769_),
    .S1(_02770_),
    .Z(_02849_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _07197_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[24][7] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[25][7] ),
    .I2(\soc.spi_video_ram_1.write_fifo.fifo_mem[26][7] ),
    .I3(\soc.spi_video_ram_1.write_fifo.fifo_mem[27][7] ),
    .S0(_02769_),
    .S1(_02770_),
    .Z(_02850_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _07198_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[20][7] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[21][7] ),
    .I2(\soc.spi_video_ram_1.write_fifo.fifo_mem[22][7] ),
    .I3(\soc.spi_video_ram_1.write_fifo.fifo_mem[23][7] ),
    .S0(_02764_),
    .S1(_02723_),
    .Z(_02851_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _07199_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[16][7] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[17][7] ),
    .I2(\soc.spi_video_ram_1.write_fifo.fifo_mem[18][7] ),
    .I3(\soc.spi_video_ram_1.write_fifo.fifo_mem[19][7] ),
    .S0(_02769_),
    .S1(_02770_),
    .Z(_02852_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _07200_ (.I0(_02849_),
    .I1(_02850_),
    .I2(_02851_),
    .I3(_02852_),
    .S0(_02571_),
    .S1(_02602_),
    .Z(_02853_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _07201_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[12][7] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[13][7] ),
    .I2(\soc.spi_video_ram_1.write_fifo.fifo_mem[14][7] ),
    .I3(\soc.spi_video_ram_1.write_fifo.fifo_mem[15][7] ),
    .S0(_02680_),
    .S1(_02838_),
    .Z(_02854_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _07202_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[8][7] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[9][7] ),
    .I2(\soc.spi_video_ram_1.write_fifo.fifo_mem[10][7] ),
    .I3(\soc.spi_video_ram_1.write_fifo.fifo_mem[11][7] ),
    .S0(_02680_),
    .S1(_02722_),
    .Z(_02855_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _07203_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[4][7] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[5][7] ),
    .I2(\soc.spi_video_ram_1.write_fifo.fifo_mem[6][7] ),
    .I3(\soc.spi_video_ram_1.write_fifo.fifo_mem[7][7] ),
    .S0(_02763_),
    .S1(_02838_),
    .Z(_02856_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _07204_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[0][7] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[1][7] ),
    .I2(\soc.spi_video_ram_1.write_fifo.fifo_mem[2][7] ),
    .I3(\soc.spi_video_ram_1.write_fifo.fifo_mem[3][7] ),
    .S0(_02680_),
    .S1(_02838_),
    .Z(_02857_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _07205_ (.I0(_02854_),
    .I1(_02855_),
    .I2(_02856_),
    .I3(_02857_),
    .S0(_02570_),
    .S1(_02719_),
    .Z(_02858_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _07206_ (.A1(_02620_),
    .A2(_02858_),
    .Z(_02859_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07207_ (.A1(_02710_),
    .A2(_02853_),
    .B(_02859_),
    .C(_02606_),
    .ZN(_02860_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07208_ (.A1(_01510_),
    .A2(_02676_),
    .B1(_02848_),
    .B2(_02860_),
    .ZN(_00240_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _07209_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[8][8] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[9][8] ),
    .I2(\soc.spi_video_ram_1.write_fifo.fifo_mem[10][8] ),
    .I3(\soc.spi_video_ram_1.write_fifo.fifo_mem[11][8] ),
    .S0(_02575_),
    .S1(_02578_),
    .Z(_02861_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07210_ (.A1(_02583_),
    .A2(_02861_),
    .ZN(_02862_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _07211_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[12][8] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[13][8] ),
    .I2(\soc.spi_video_ram_1.write_fifo.fifo_mem[14][8] ),
    .I3(\soc.spi_video_ram_1.write_fifo.fifo_mem[15][8] ),
    .S0(_02575_),
    .S1(_02578_),
    .Z(_02863_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07212_ (.A1(_02571_),
    .A2(_02863_),
    .B(_02586_),
    .ZN(_02864_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _07213_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[0][8] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[1][8] ),
    .I2(\soc.spi_video_ram_1.write_fifo.fifo_mem[2][8] ),
    .I3(\soc.spi_video_ram_1.write_fifo.fifo_mem[3][8] ),
    .S0(_02591_),
    .S1(_02593_),
    .Z(_02865_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07214_ (.A1(_02589_),
    .A2(_02865_),
    .ZN(_02866_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _07215_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[4][8] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[5][8] ),
    .I2(\soc.spi_video_ram_1.write_fifo.fifo_mem[6][8] ),
    .I3(\soc.spi_video_ram_1.write_fifo.fifo_mem[7][8] ),
    .S0(_02597_),
    .S1(_02598_),
    .Z(_02867_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07216_ (.A1(_02596_),
    .A2(_02867_),
    .B(_02618_),
    .ZN(_02868_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _07217_ (.A1(_02862_),
    .A2(_02864_),
    .B1(_02866_),
    .B2(_02868_),
    .ZN(_02869_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07218_ (.A1(_02568_),
    .A2(_02869_),
    .ZN(_02870_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _07219_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[28][8] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[29][8] ),
    .I2(\soc.spi_video_ram_1.write_fifo.fifo_mem[30][8] ),
    .I3(\soc.spi_video_ram_1.write_fifo.fifo_mem[31][8] ),
    .S0(_02607_),
    .S1(_02636_),
    .Z(_02871_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07220_ (.A1(_02596_),
    .A2(_02871_),
    .ZN(_02872_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _07221_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[24][8] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[25][8] ),
    .I2(\soc.spi_video_ram_1.write_fifo.fifo_mem[26][8] ),
    .I3(\soc.spi_video_ram_1.write_fifo.fifo_mem[27][8] ),
    .S0(_02607_),
    .S1(_02578_),
    .Z(_02873_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07222_ (.A1(_02583_),
    .A2(_02873_),
    .B(_02640_),
    .ZN(_02874_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _07223_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[16][8] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[17][8] ),
    .I2(\soc.spi_video_ram_1.write_fifo.fifo_mem[18][8] ),
    .I3(\soc.spi_video_ram_1.write_fifo.fifo_mem[19][8] ),
    .S0(_02645_),
    .S1(_02614_),
    .Z(_02875_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07224_ (.A1(_02589_),
    .A2(_02875_),
    .ZN(_02876_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _07225_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[20][8] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[21][8] ),
    .I2(\soc.spi_video_ram_1.write_fifo.fifo_mem[22][8] ),
    .I3(\soc.spi_video_ram_1.write_fifo.fifo_mem[23][8] ),
    .S0(_02591_),
    .S1(_02593_),
    .Z(_02877_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07226_ (.A1(_02650_),
    .A2(_02877_),
    .B(_02618_),
    .ZN(_02878_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _07227_ (.A1(_02872_),
    .A2(_02874_),
    .B1(_02876_),
    .B2(_02878_),
    .C(_02620_),
    .ZN(_02879_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07228_ (.A1(_02606_),
    .A2(_02879_),
    .ZN(_02880_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07229_ (.A1(_02870_),
    .A2(_02880_),
    .B(_02626_),
    .ZN(_02881_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07230_ (.I(_02734_),
    .Z(_02882_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07231_ (.I0(\soc.spi_video_ram_1.output_buffer[15] ),
    .I1(_02881_),
    .S(_02882_),
    .Z(_02883_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07232_ (.I(_02883_),
    .Z(_00241_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _07233_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[12][9] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[13][9] ),
    .I2(\soc.spi_video_ram_1.write_fifo.fifo_mem[14][9] ),
    .I3(\soc.spi_video_ram_1.write_fifo.fifo_mem[15][9] ),
    .S0(_02645_),
    .S1(_02614_),
    .Z(_02884_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07234_ (.A1(_02650_),
    .A2(_02884_),
    .ZN(_02885_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _07235_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[8][9] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[9][9] ),
    .I2(\soc.spi_video_ram_1.write_fifo.fifo_mem[10][9] ),
    .I3(\soc.spi_video_ram_1.write_fifo.fifo_mem[11][9] ),
    .S0(_02645_),
    .S1(_02614_),
    .Z(_02886_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07236_ (.A1(_02589_),
    .A2(_02886_),
    .B(_02640_),
    .ZN(_02887_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _07237_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[0][9] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[1][9] ),
    .I2(\soc.spi_video_ram_1.write_fifo.fifo_mem[2][9] ),
    .I3(\soc.spi_video_ram_1.write_fifo.fifo_mem[3][9] ),
    .S0(_02680_),
    .S1(_02722_),
    .Z(_02888_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07238_ (.A1(_02643_),
    .A2(_02888_),
    .ZN(_02889_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _07239_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[4][9] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[5][9] ),
    .I2(\soc.spi_video_ram_1.write_fifo.fifo_mem[6][9] ),
    .I3(\soc.spi_video_ram_1.write_fifo.fifo_mem[7][9] ),
    .S0(_02712_),
    .S1(_02722_),
    .Z(_02890_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07240_ (.A1(_02650_),
    .A2(_02890_),
    .B(_02719_),
    .ZN(_02891_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _07241_ (.A1(_02885_),
    .A2(_02887_),
    .B1(_02889_),
    .B2(_02891_),
    .ZN(_02892_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 _07242_ (.I(_02679_),
    .Z(_02893_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07243_ (.I(_02576_),
    .Z(_02894_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07244_ (.I(_02894_),
    .Z(_02895_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _07245_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[28][9] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[29][9] ),
    .I2(\soc.spi_video_ram_1.write_fifo.fifo_mem[30][9] ),
    .I3(\soc.spi_video_ram_1.write_fifo.fifo_mem[31][9] ),
    .S0(_02893_),
    .S1(_02895_),
    .Z(_02896_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07246_ (.A1(_02570_),
    .A2(_02896_),
    .ZN(_02897_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _07247_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[24][9] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[25][9] ),
    .I2(\soc.spi_video_ram_1.write_fifo.fifo_mem[26][9] ),
    .I3(\soc.spi_video_ram_1.write_fifo.fifo_mem[27][9] ),
    .S0(_02893_),
    .S1(_02827_),
    .Z(_02898_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07248_ (.A1(_02767_),
    .A2(_02898_),
    .B(_02831_),
    .ZN(_02899_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07249_ (.I(_00002_),
    .Z(_02900_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07250_ (.I(_02900_),
    .Z(_02901_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _07251_ (.I(_02572_),
    .Z(_02902_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 _07252_ (.I(_02902_),
    .Z(_02903_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _07253_ (.I(_02894_),
    .Z(_02904_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _07254_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[16][9] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[17][9] ),
    .I2(\soc.spi_video_ram_1.write_fifo.fifo_mem[18][9] ),
    .I3(\soc.spi_video_ram_1.write_fifo.fifo_mem[19][9] ),
    .S0(_02903_),
    .S1(_02904_),
    .Z(_02905_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07255_ (.A1(_02901_),
    .A2(_02905_),
    .ZN(_02906_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 _07256_ (.I(_02679_),
    .Z(_02907_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07257_ (.I(_02894_),
    .Z(_02908_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _07258_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[20][9] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[21][9] ),
    .I2(\soc.spi_video_ram_1.write_fifo.fifo_mem[22][9] ),
    .I3(\soc.spi_video_ram_1.write_fifo.fifo_mem[23][9] ),
    .S0(_02907_),
    .S1(_02908_),
    .Z(_02909_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07259_ (.I(_02600_),
    .Z(_02910_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07260_ (.A1(_02570_),
    .A2(_02909_),
    .B(_02910_),
    .ZN(_02911_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _07261_ (.A1(_02897_),
    .A2(_02899_),
    .B1(_02906_),
    .B2(_02911_),
    .C(_02567_),
    .ZN(_02912_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07262_ (.A1(_02620_),
    .A2(_02892_),
    .B(_02912_),
    .C(_02606_),
    .ZN(_02913_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07263_ (.A1(_02058_),
    .A2(_02625_),
    .B(_02913_),
    .ZN(_02914_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07264_ (.I0(\soc.spi_video_ram_1.output_buffer[14] ),
    .I1(_02914_),
    .S(_02633_),
    .Z(_02915_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07265_ (.I(_02915_),
    .Z(_00242_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07266_ (.I(_02056_),
    .ZN(_02916_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07267_ (.A1(_02055_),
    .A2(_02916_),
    .Z(_02917_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _07268_ (.A1(_01387_),
    .A2(_01386_),
    .A3(\soc.spi_video_ram_1.state_sram_clk_counter[0] ),
    .A4(_01390_),
    .ZN(_02918_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _07269_ (.I(_02573_),
    .Z(_02919_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07270_ (.I(_02919_),
    .Z(_02920_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07271_ (.A1(_02920_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[10][10] ),
    .ZN(_02921_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07272_ (.I(_02695_),
    .Z(_02922_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07273_ (.A1(_02922_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[11][10] ),
    .B(_02647_),
    .ZN(_02923_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07274_ (.I(_02590_),
    .Z(_02924_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07275_ (.A1(_02924_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[8][10] ),
    .ZN(_02925_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07276_ (.I(_02695_),
    .Z(_02926_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07277_ (.I(_02740_),
    .Z(_02927_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07278_ (.A1(_02926_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[9][10] ),
    .B(_02927_),
    .ZN(_02928_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07279_ (.I(_02569_),
    .Z(_02929_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _07280_ (.A1(_02921_),
    .A2(_02923_),
    .B1(_02925_),
    .B2(_02928_),
    .C(_02929_),
    .ZN(_02930_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07281_ (.I(_02573_),
    .Z(_02931_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _07282_ (.A1(_02931_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[13][10] ),
    .Z(_02932_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07283_ (.A1(_02922_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[12][10] ),
    .B(_02932_),
    .ZN(_02933_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07284_ (.A1(_02924_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[14][10] ),
    .ZN(_02934_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07285_ (.A1(_02926_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[15][10] ),
    .B(_02838_),
    .ZN(_02935_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _07286_ (.A1(_02691_),
    .A2(_02933_),
    .B1(_02934_),
    .B2(_02935_),
    .C(_02588_),
    .ZN(_02936_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07287_ (.A1(_02831_),
    .A2(_02930_),
    .A3(_02936_),
    .ZN(_02937_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _07288_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[0][10] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[1][10] ),
    .I2(\soc.spi_video_ram_1.write_fifo.fifo_mem[2][10] ),
    .I3(\soc.spi_video_ram_1.write_fifo.fifo_mem[3][10] ),
    .S0(_02893_),
    .S1(_02895_),
    .Z(_02938_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07289_ (.A1(_02696_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[7][10] ),
    .ZN(_02939_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07290_ (.A1(_02744_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[6][10] ),
    .B(_02895_),
    .ZN(_02940_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07291_ (.I(_02694_),
    .Z(_02941_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07292_ (.A1(_02941_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[5][10] ),
    .ZN(_02942_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07293_ (.I(_02740_),
    .Z(_02943_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07294_ (.A1(_02597_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[4][10] ),
    .B(_02943_),
    .ZN(_02944_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _07295_ (.A1(_02939_),
    .A2(_02940_),
    .B1(_02942_),
    .B2(_02944_),
    .C(_02706_),
    .ZN(_02945_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07296_ (.A1(_02707_),
    .A2(_02938_),
    .B(_02945_),
    .C(_02910_),
    .ZN(_02946_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07297_ (.A1(_02937_),
    .A2(_02946_),
    .ZN(_02947_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07298_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[18][10] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[19][10] ),
    .S(_02893_),
    .Z(_02948_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07299_ (.A1(_02597_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[17][10] ),
    .ZN(_02949_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07300_ (.A1(_02941_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[16][10] ),
    .ZN(_02950_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07301_ (.A1(_02949_),
    .A2(_02950_),
    .B(_02598_),
    .ZN(_02951_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07302_ (.I(_02581_),
    .Z(_02952_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _07303_ (.A1(_02758_),
    .A2(_02948_),
    .B(_02951_),
    .C(_02952_),
    .ZN(_02953_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07304_ (.A1(_02744_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[22][10] ),
    .ZN(_02954_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07305_ (.A1(_02696_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[23][10] ),
    .B(_02895_),
    .ZN(_02955_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _07306_ (.A1(_02612_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[21][10] ),
    .Z(_02956_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07307_ (.A1(_02941_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[20][10] ),
    .B(_02956_),
    .ZN(_02957_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07308_ (.I(_02577_),
    .Z(_02958_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _07309_ (.A1(_02954_),
    .A2(_02955_),
    .B1(_02957_),
    .B2(_02958_),
    .C(_02642_),
    .ZN(_02959_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07310_ (.A1(_02910_),
    .A2(_02959_),
    .ZN(_02960_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _07311_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[24][10] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[25][10] ),
    .I2(\soc.spi_video_ram_1.write_fifo.fifo_mem[26][10] ),
    .I3(\soc.spi_video_ram_1.write_fifo.fifo_mem[27][10] ),
    .S0(_02574_),
    .S1(_02592_),
    .Z(_02961_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07312_ (.A1(_02703_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[31][10] ),
    .ZN(_02962_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07313_ (.A1(_02763_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[30][10] ),
    .B(_02592_),
    .ZN(_02963_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _07314_ (.A1(_02573_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[29][10] ),
    .Z(_02964_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07315_ (.A1(_02703_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[28][10] ),
    .B(_02964_),
    .ZN(_02965_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _07316_ (.A1(_02962_),
    .A2(_02963_),
    .B1(_02965_),
    .B2(_02722_),
    .C(_02900_),
    .ZN(_02966_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07317_ (.A1(_02952_),
    .A2(_02961_),
    .B(_02966_),
    .C(_02585_),
    .ZN(_02967_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07318_ (.A1(_02953_),
    .A2(_02960_),
    .B(_00004_),
    .C(_02967_),
    .ZN(_02968_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07319_ (.A1(_02620_),
    .A2(_02947_),
    .B(_02968_),
    .ZN(_02969_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07320_ (.I(_00003_),
    .Z(_02970_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07321_ (.I(_02574_),
    .Z(_02971_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07322_ (.A1(_02971_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[14][28] ),
    .ZN(_02972_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07323_ (.A1(_02926_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[15][28] ),
    .B(_02722_),
    .ZN(_02973_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _07324_ (.A1(_02590_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[13][28] ),
    .Z(_02974_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07325_ (.A1(_02696_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[12][28] ),
    .B(_02974_),
    .ZN(_02975_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07326_ (.I(_02577_),
    .Z(_02976_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _07327_ (.A1(_02972_),
    .A2(_02973_),
    .B1(_02975_),
    .B2(_02976_),
    .C(_02642_),
    .ZN(_02977_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07328_ (.A1(_02971_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[10][28] ),
    .ZN(_02978_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07329_ (.A1(_02922_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[11][28] ),
    .B(_02722_),
    .ZN(_02979_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07330_ (.A1(_02744_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[8][28] ),
    .ZN(_02980_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07331_ (.A1(_02696_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[9][28] ),
    .B(_02927_),
    .ZN(_02981_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _07332_ (.A1(_02978_),
    .A2(_02979_),
    .B1(_02980_),
    .B2(_02981_),
    .C(_02569_),
    .ZN(_02982_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _07333_ (.A1(_02970_),
    .A2(_02977_),
    .A3(_02982_),
    .Z(_02983_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07334_ (.I(_02900_),
    .Z(_02984_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _07335_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[0][28] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[1][28] ),
    .I2(\soc.spi_video_ram_1.write_fifo.fifo_mem[2][28] ),
    .I3(\soc.spi_video_ram_1.write_fifo.fifo_mem[3][28] ),
    .S0(_02931_),
    .S1(_02690_),
    .Z(_02985_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07336_ (.A1(_02941_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[7][28] ),
    .ZN(_02986_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07337_ (.A1(_02651_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[6][28] ),
    .B(_02690_),
    .ZN(_02987_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07338_ (.A1(_02703_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[5][28] ),
    .ZN(_02988_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07339_ (.A1(_02712_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[4][28] ),
    .B(_02741_),
    .ZN(_02989_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _07340_ (.A1(_02986_),
    .A2(_02987_),
    .B1(_02988_),
    .B2(_02989_),
    .C(_02900_),
    .ZN(_02990_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07341_ (.A1(_02984_),
    .A2(_02985_),
    .B(_02990_),
    .C(_02601_),
    .ZN(_02991_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07342_ (.A1(_02655_),
    .A2(_02991_),
    .ZN(_02992_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07343_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[18][28] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[19][28] ),
    .S(_02783_),
    .Z(_02993_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07344_ (.A1(_02712_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[17][28] ),
    .ZN(_02994_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07345_ (.A1(_02703_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[16][28] ),
    .ZN(_02995_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07346_ (.A1(_02994_),
    .A2(_02995_),
    .B(_02838_),
    .ZN(_02996_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _07347_ (.A1(_02691_),
    .A2(_02993_),
    .B(_02996_),
    .C(_02582_),
    .ZN(_02997_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07348_ (.A1(_02613_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[22][28] ),
    .ZN(_02998_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07349_ (.A1(_02941_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[23][28] ),
    .B(_02690_),
    .ZN(_02999_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _07350_ (.A1(_02679_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[21][28] ),
    .Z(_03000_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07351_ (.A1(_02703_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[20][28] ),
    .B(_03000_),
    .ZN(_03001_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _07352_ (.A1(_02998_),
    .A2(_02999_),
    .B1(_03001_),
    .B2(_02598_),
    .C(_02900_),
    .ZN(_03002_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07353_ (.A1(_02601_),
    .A2(_03002_),
    .ZN(_03003_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _07354_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[24][28] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[25][28] ),
    .I2(\soc.spi_video_ram_1.write_fifo.fifo_mem[26][28] ),
    .I3(\soc.spi_video_ram_1.write_fifo.fifo_mem[27][28] ),
    .S0(_02644_),
    .S1(_02646_),
    .Z(_03004_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07355_ (.A1(_02695_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[31][28] ),
    .ZN(_03005_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07356_ (.A1(_02903_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[30][28] ),
    .B(_02646_),
    .ZN(_03006_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _07357_ (.A1(_02573_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[29][28] ),
    .Z(_03007_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07358_ (.A1(_02695_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[28][28] ),
    .B(_03007_),
    .ZN(_03008_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _07359_ (.A1(_03005_),
    .A2(_03006_),
    .B1(_03008_),
    .B2(_02908_),
    .C(_02581_),
    .ZN(_03009_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07360_ (.A1(_02582_),
    .A2(_03004_),
    .B(_03009_),
    .C(_02585_),
    .ZN(_03010_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07361_ (.A1(_02997_),
    .A2(_03003_),
    .B(_00004_),
    .C(_03010_),
    .ZN(_03011_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07362_ (.A1(_02983_),
    .A2(_02992_),
    .B(_03011_),
    .C(_02918_),
    .ZN(_03012_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07363_ (.A1(_02918_),
    .A2(_02969_),
    .B(_03012_),
    .ZN(_03013_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07364_ (.A1(_01419_),
    .A2(_02917_),
    .B1(_03013_),
    .B2(_02677_),
    .ZN(_03014_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07365_ (.A1(_02624_),
    .A2(_02882_),
    .ZN(_03015_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07366_ (.A1(\soc.spi_video_ram_1.output_buffer[13] ),
    .A2(_02676_),
    .ZN(_03016_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07367_ (.A1(_03014_),
    .A2(_03015_),
    .B(_03016_),
    .ZN(_00243_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07368_ (.A1(_01939_),
    .A2(_02034_),
    .ZN(_03017_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07369_ (.A1(_01964_),
    .A2(_03017_),
    .B(_02916_),
    .ZN(_03018_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07370_ (.I(_02918_),
    .ZN(_03019_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07371_ (.A1(_02784_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[18][11] ),
    .ZN(_03020_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07372_ (.I(_02695_),
    .Z(_03021_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07373_ (.A1(_03021_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[19][11] ),
    .B(_02614_),
    .ZN(_03022_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07374_ (.A1(_02971_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[16][11] ),
    .ZN(_03023_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07375_ (.I(_02741_),
    .Z(_03024_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07376_ (.A1(_02922_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[17][11] ),
    .B(_03024_),
    .ZN(_03025_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _07377_ (.A1(_03020_),
    .A2(_03022_),
    .B1(_03023_),
    .B2(_03025_),
    .C(_02929_),
    .ZN(_03026_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07378_ (.A1(_02784_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[22][11] ),
    .ZN(_03027_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07379_ (.A1(_03021_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[23][11] ),
    .B(_02614_),
    .ZN(_03028_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _07380_ (.A1(_02919_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[21][11] ),
    .Z(_03029_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07381_ (.A1(_02926_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[20][11] ),
    .B(_03029_),
    .ZN(_03030_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _07382_ (.A1(_03027_),
    .A2(_03028_),
    .B1(_03030_),
    .B2(_02691_),
    .C(_02588_),
    .ZN(_03031_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07383_ (.A1(_02719_),
    .A2(_03026_),
    .A3(_03031_),
    .ZN(_03032_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _07384_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[24][11] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[25][11] ),
    .I2(\soc.spi_video_ram_1.write_fifo.fifo_mem[26][11] ),
    .I3(\soc.spi_video_ram_1.write_fifo.fifo_mem[27][11] ),
    .S0(_02688_),
    .S1(_02827_),
    .Z(_03033_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07385_ (.A1(_02696_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[31][11] ),
    .ZN(_03034_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07386_ (.A1(_02924_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[30][11] ),
    .B(_02827_),
    .ZN(_03035_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _07387_ (.A1(_02612_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[29][11] ),
    .Z(_03036_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07388_ (.A1(_02696_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[28][11] ),
    .B(_03036_),
    .ZN(_03037_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _07389_ (.A1(_03034_),
    .A2(_03035_),
    .B1(_03037_),
    .B2(_02976_),
    .C(_02642_),
    .ZN(_03038_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07390_ (.A1(_02767_),
    .A2(_03033_),
    .B(_03038_),
    .C(_02831_),
    .ZN(_03039_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07391_ (.A1(_02620_),
    .A2(_03032_),
    .A3(_03039_),
    .ZN(_03040_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07392_ (.I(_02958_),
    .Z(_03041_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07393_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[14][11] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[15][11] ),
    .S(_02613_),
    .Z(_03042_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07394_ (.A1(_02920_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[13][11] ),
    .ZN(_03043_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07395_ (.A1(_02926_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[12][11] ),
    .ZN(_03044_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07396_ (.A1(_03043_),
    .A2(_03044_),
    .B(_02958_),
    .ZN(_03045_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _07397_ (.A1(_03041_),
    .A2(_03042_),
    .B(_03045_),
    .C(_02570_),
    .ZN(_03046_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07398_ (.I(_02783_),
    .Z(_03047_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07399_ (.A1(_03047_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[10][11] ),
    .ZN(_03048_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07400_ (.A1(_03021_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[11][11] ),
    .B(_02652_),
    .ZN(_03049_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07401_ (.A1(_02971_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[8][11] ),
    .ZN(_03050_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07402_ (.A1(_02922_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[9][11] ),
    .B(_03024_),
    .ZN(_03051_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _07403_ (.A1(_03048_),
    .A2(_03049_),
    .B1(_03050_),
    .B2(_03051_),
    .C(_02929_),
    .ZN(_03052_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07404_ (.A1(_02640_),
    .A2(_03052_),
    .ZN(_03053_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 _07405_ (.I(_02902_),
    .Z(_03054_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _07406_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[0][11] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[1][11] ),
    .I2(\soc.spi_video_ram_1.write_fifo.fifo_mem[2][11] ),
    .I3(\soc.spi_video_ram_1.write_fifo.fifo_mem[3][11] ),
    .S0(_03054_),
    .S1(_02690_),
    .Z(_03055_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _07407_ (.A1(_02644_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[4][11] ),
    .Z(_03056_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07408_ (.A1(_02941_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[5][11] ),
    .B(_03056_),
    .ZN(_03057_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07409_ (.A1(_02941_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[7][11] ),
    .ZN(_03058_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07410_ (.A1(_02700_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[6][11] ),
    .B(_02577_),
    .ZN(_03059_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _07411_ (.A1(_02578_),
    .A2(_03057_),
    .B1(_03058_),
    .B2(_03059_),
    .C(_02900_),
    .ZN(_03060_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07412_ (.A1(_02901_),
    .A2(_03055_),
    .B(_03060_),
    .C(_02910_),
    .ZN(_03061_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07413_ (.A1(_03046_),
    .A2(_03053_),
    .B(_03061_),
    .C(_02655_),
    .ZN(_03062_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07414_ (.A1(_03019_),
    .A2(_03040_),
    .A3(_03062_),
    .ZN(_03063_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07415_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[14][27] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[15][27] ),
    .S(_02613_),
    .Z(_03064_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07416_ (.A1(_02971_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[13][27] ),
    .ZN(_03065_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07417_ (.A1(_02696_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[12][27] ),
    .ZN(_03066_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07418_ (.A1(_03065_),
    .A2(_03066_),
    .B(_02958_),
    .ZN(_03067_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _07419_ (.A1(_03041_),
    .A2(_03064_),
    .B(_03067_),
    .C(_02570_),
    .ZN(_03068_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07420_ (.A1(_02784_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[10][27] ),
    .ZN(_03069_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07421_ (.A1(_03021_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[11][27] ),
    .B(_02652_),
    .ZN(_03070_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07422_ (.A1(_02971_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[8][27] ),
    .ZN(_03071_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07423_ (.A1(_02922_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[9][27] ),
    .B(_03024_),
    .ZN(_03072_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _07424_ (.A1(_03069_),
    .A2(_03070_),
    .B1(_03071_),
    .B2(_03072_),
    .C(_02929_),
    .ZN(_03073_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07425_ (.A1(_02831_),
    .A2(_03073_),
    .ZN(_03074_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _07426_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[0][27] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[1][27] ),
    .I2(\soc.spi_video_ram_1.write_fifo.fifo_mem[2][27] ),
    .I3(\soc.spi_video_ram_1.write_fifo.fifo_mem[3][27] ),
    .S0(_03054_),
    .S1(_02690_),
    .Z(_03075_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07427_ (.A1(_02941_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[7][27] ),
    .ZN(_03076_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07428_ (.A1(_02597_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[6][27] ),
    .B(_02690_),
    .ZN(_03077_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07429_ (.A1(_02703_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[5][27] ),
    .ZN(_03078_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07430_ (.A1(_02700_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[4][27] ),
    .B(_02943_),
    .ZN(_03079_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _07431_ (.A1(_03076_),
    .A2(_03077_),
    .B1(_03078_),
    .B2(_03079_),
    .C(_02900_),
    .ZN(_03080_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07432_ (.A1(_02901_),
    .A2(_03075_),
    .B(_03080_),
    .C(_02910_),
    .ZN(_03081_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07433_ (.A1(_03068_),
    .A2(_03074_),
    .B(_03081_),
    .C(_02655_),
    .ZN(_03082_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _07434_ (.A1(_03054_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[21][27] ),
    .Z(_03083_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07435_ (.A1(_03021_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[20][27] ),
    .B(_03083_),
    .ZN(_03084_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07436_ (.A1(_02752_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[22][27] ),
    .ZN(_03085_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07437_ (.A1(_02922_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[23][27] ),
    .B(_02722_),
    .ZN(_03086_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _07438_ (.A1(_02691_),
    .A2(_03084_),
    .B1(_03085_),
    .B2(_03086_),
    .C(_02588_),
    .ZN(_03087_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07439_ (.A1(_02784_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[18][27] ),
    .ZN(_03088_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07440_ (.A1(_03021_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[19][27] ),
    .B(_02614_),
    .ZN(_03089_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07441_ (.A1(_02752_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[16][27] ),
    .ZN(_03090_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07442_ (.A1(_02926_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[17][27] ),
    .B(_03024_),
    .ZN(_03091_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _07443_ (.A1(_03088_),
    .A2(_03089_),
    .B1(_03090_),
    .B2(_03091_),
    .C(_02929_),
    .ZN(_03092_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07444_ (.A1(_02719_),
    .A2(_03087_),
    .A3(_03092_),
    .ZN(_03093_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _07445_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[24][27] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[25][27] ),
    .I2(\soc.spi_video_ram_1.write_fifo.fifo_mem[26][27] ),
    .I3(\soc.spi_video_ram_1.write_fifo.fifo_mem[27][27] ),
    .S0(_02688_),
    .S1(_02827_),
    .Z(_03094_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07446_ (.A1(_02696_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[31][27] ),
    .ZN(_03095_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07447_ (.A1(_02924_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[30][27] ),
    .B(_02827_),
    .ZN(_03096_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _07448_ (.A1(_02612_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[29][27] ),
    .Z(_03097_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07449_ (.A1(_02696_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[28][27] ),
    .B(_03097_),
    .ZN(_03098_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _07450_ (.A1(_03095_),
    .A2(_03096_),
    .B1(_03098_),
    .B2(_02958_),
    .C(_02642_),
    .ZN(_03099_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07451_ (.A1(_02767_),
    .A2(_03094_),
    .B(_03099_),
    .C(_02970_),
    .ZN(_03100_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07452_ (.A1(_02567_),
    .A2(_03093_),
    .A3(_03100_),
    .ZN(_03101_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07453_ (.A1(_02918_),
    .A2(_03082_),
    .A3(_03101_),
    .ZN(_03102_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07454_ (.A1(_03063_),
    .A2(_03102_),
    .ZN(_03103_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07455_ (.A1(_01419_),
    .A2(_03018_),
    .B1(_03103_),
    .B2(_02677_),
    .ZN(_03104_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07456_ (.A1(\soc.spi_video_ram_1.output_buffer[12] ),
    .A2(_02676_),
    .ZN(_03105_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07457_ (.A1(_03015_),
    .A2(_03104_),
    .B(_03105_),
    .ZN(_00244_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07458_ (.A1(_01939_),
    .A2(_01930_),
    .Z(_03106_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07459_ (.A1(_01940_),
    .A2(_03106_),
    .ZN(_03107_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _07460_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[16][12] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[17][12] ),
    .I2(\soc.spi_video_ram_1.write_fifo.fifo_mem[18][12] ),
    .I3(\soc.spi_video_ram_1.write_fifo.fifo_mem[19][12] ),
    .S0(_02903_),
    .S1(_02904_),
    .Z(_03108_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07461_ (.I(\soc.spi_video_ram_1.write_fifo.fifo_mem[23][12] ),
    .ZN(_03109_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07462_ (.A1(_03054_),
    .A2(_03109_),
    .ZN(_03110_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07463_ (.A1(_02607_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[22][12] ),
    .B(_03110_),
    .C(_02904_),
    .ZN(_03111_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07464_ (.I(\soc.spi_video_ram_1.write_fifo.fifo_mem[21][12] ),
    .ZN(_03112_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07465_ (.A1(_03054_),
    .A2(_03112_),
    .ZN(_03113_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07466_ (.A1(_02607_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[20][12] ),
    .B(_03113_),
    .C(_02943_),
    .ZN(_03114_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07467_ (.A1(_02642_),
    .A2(_03111_),
    .A3(_03114_),
    .ZN(_03115_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07468_ (.A1(_02901_),
    .A2(_03108_),
    .B(_03115_),
    .C(_02910_),
    .ZN(_03116_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _07469_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[24][12] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[25][12] ),
    .I2(\soc.spi_video_ram_1.write_fifo.fifo_mem[26][12] ),
    .I3(\soc.spi_video_ram_1.write_fifo.fifo_mem[27][12] ),
    .S0(_03054_),
    .S1(_02904_),
    .Z(_03117_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07470_ (.I(\soc.spi_video_ram_1.write_fifo.fifo_mem[29][12] ),
    .ZN(_03118_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07471_ (.A1(_02931_),
    .A2(_03118_),
    .ZN(_03119_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07472_ (.A1(_02597_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[28][12] ),
    .B(_03119_),
    .C(_02943_),
    .ZN(_03120_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07473_ (.I(\soc.spi_video_ram_1.write_fifo.fifo_mem[31][12] ),
    .ZN(_03121_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07474_ (.A1(_02931_),
    .A2(_03121_),
    .ZN(_03122_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07475_ (.A1(_02597_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[30][12] ),
    .B(_03122_),
    .C(_02904_),
    .ZN(_03123_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07476_ (.A1(_02642_),
    .A2(_03120_),
    .A3(_03123_),
    .ZN(_03124_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07477_ (.A1(_02901_),
    .A2(_03117_),
    .B(_03124_),
    .C(_02970_),
    .ZN(_03125_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07478_ (.A1(_03116_),
    .A2(_03125_),
    .ZN(_03126_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _07479_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[0][12] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[1][12] ),
    .I2(\soc.spi_video_ram_1.write_fifo.fifo_mem[2][12] ),
    .I3(\soc.spi_video_ram_1.write_fifo.fifo_mem[3][12] ),
    .S0(_02919_),
    .S1(_02577_),
    .Z(_03127_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07480_ (.I(\soc.spi_video_ram_1.write_fifo.fifo_mem[5][12] ),
    .ZN(_03128_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07481_ (.A1(_02919_),
    .A2(_03128_),
    .ZN(_03129_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07482_ (.A1(_02613_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[4][12] ),
    .B(_03129_),
    .C(_02943_),
    .ZN(_03130_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07483_ (.I(\soc.spi_video_ram_1.write_fifo.fifo_mem[7][12] ),
    .ZN(_03131_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07484_ (.A1(_02919_),
    .A2(_03131_),
    .ZN(_03132_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07485_ (.A1(_02645_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[6][12] ),
    .B(_03132_),
    .C(_02577_),
    .ZN(_03133_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07486_ (.A1(_02706_),
    .A2(_03130_),
    .A3(_03133_),
    .ZN(_03134_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07487_ (.A1(_02984_),
    .A2(_03127_),
    .B(_03134_),
    .C(_02601_),
    .ZN(_03135_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _07488_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[8][12] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[9][12] ),
    .I2(\soc.spi_video_ram_1.write_fifo.fifo_mem[10][12] ),
    .I3(\soc.spi_video_ram_1.write_fifo.fifo_mem[11][12] ),
    .S0(_02574_),
    .S1(_02577_),
    .Z(_03136_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07489_ (.A1(_02941_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[13][12] ),
    .ZN(_03137_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07490_ (.A1(_02712_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[12][12] ),
    .B(_02943_),
    .ZN(_03138_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _07491_ (.I(_02679_),
    .Z(_03139_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07492_ (.I(\soc.spi_video_ram_1.write_fifo.fifo_mem[15][12] ),
    .ZN(_03140_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07493_ (.A1(_02644_),
    .A2(_03140_),
    .ZN(_03141_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07494_ (.A1(_03139_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[14][12] ),
    .B(_03141_),
    .C(_02646_),
    .ZN(_03142_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07495_ (.A1(_03137_),
    .A2(_03138_),
    .B(_02900_),
    .C(_03142_),
    .ZN(_03143_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07496_ (.A1(_02952_),
    .A2(_03136_),
    .B(_03143_),
    .C(_02585_),
    .ZN(_03144_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07497_ (.A1(_03135_),
    .A2(_03144_),
    .B(_02567_),
    .ZN(_03145_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _07498_ (.A1(_02620_),
    .A2(_03126_),
    .B(_03145_),
    .C(_02918_),
    .ZN(_03146_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _07499_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[16][26] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[17][26] ),
    .I2(\soc.spi_video_ram_1.write_fifo.fifo_mem[18][26] ),
    .I3(\soc.spi_video_ram_1.write_fifo.fifo_mem[19][26] ),
    .S0(_02907_),
    .S1(_02908_),
    .Z(_03147_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07500_ (.I(\soc.spi_video_ram_1.write_fifo.fifo_mem[21][26] ),
    .ZN(_03148_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07501_ (.A1(_02903_),
    .A2(_03148_),
    .ZN(_03149_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07502_ (.A1(_02744_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[20][26] ),
    .B(_03149_),
    .C(_02927_),
    .ZN(_03150_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07503_ (.I(\soc.spi_video_ram_1.write_fifo.fifo_mem[23][26] ),
    .ZN(_03151_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07504_ (.A1(_02903_),
    .A2(_03151_),
    .ZN(_03152_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07505_ (.A1(_02744_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[22][26] ),
    .B(_03152_),
    .C(_02908_),
    .ZN(_03153_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07506_ (.A1(_02588_),
    .A2(_03150_),
    .A3(_03153_),
    .ZN(_03154_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07507_ (.A1(_02707_),
    .A2(_03147_),
    .B(_03154_),
    .C(_02910_),
    .ZN(_03155_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _07508_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[24][26] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[25][26] ),
    .I2(\soc.spi_video_ram_1.write_fifo.fifo_mem[26][26] ),
    .I3(\soc.spi_video_ram_1.write_fifo.fifo_mem[27][26] ),
    .S0(_02907_),
    .S1(_02908_),
    .Z(_03156_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07509_ (.I(\soc.spi_video_ram_1.write_fifo.fifo_mem[31][26] ),
    .ZN(_03157_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07510_ (.A1(_02903_),
    .A2(_03157_),
    .ZN(_03158_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07511_ (.A1(_02744_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[30][26] ),
    .B(_03158_),
    .C(_02908_),
    .ZN(_03159_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07512_ (.I(\soc.spi_video_ram_1.write_fifo.fifo_mem[29][26] ),
    .ZN(_03160_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07513_ (.A1(_02903_),
    .A2(_03160_),
    .ZN(_03161_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07514_ (.A1(_02575_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[28][26] ),
    .B(_03161_),
    .C(_02927_),
    .ZN(_03162_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07515_ (.A1(_02588_),
    .A2(_03159_),
    .A3(_03162_),
    .ZN(_03163_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07516_ (.A1(_02707_),
    .A2(_03156_),
    .B(_03163_),
    .C(_02970_),
    .ZN(_03164_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07517_ (.A1(_03155_),
    .A2(_03164_),
    .ZN(_03165_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _07518_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[8][26] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[9][26] ),
    .I2(\soc.spi_video_ram_1.write_fifo.fifo_mem[10][26] ),
    .I3(\soc.spi_video_ram_1.write_fifo.fifo_mem[11][26] ),
    .S0(_02783_),
    .S1(_02690_),
    .Z(_03166_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07519_ (.A1(_02941_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[13][26] ),
    .ZN(_03167_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07520_ (.A1(_02597_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[12][26] ),
    .B(_02943_),
    .ZN(_03168_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07521_ (.I(\soc.spi_video_ram_1.write_fifo.fifo_mem[15][26] ),
    .ZN(_03169_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07522_ (.A1(_02590_),
    .A2(_03169_),
    .ZN(_03170_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07523_ (.A1(_02763_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[14][26] ),
    .B(_03170_),
    .C(_02592_),
    .ZN(_03171_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07524_ (.A1(_03167_),
    .A2(_03168_),
    .B(_03171_),
    .C(_02706_),
    .ZN(_03172_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07525_ (.A1(_02984_),
    .A2(_03166_),
    .B(_03172_),
    .C(_02585_),
    .ZN(_03173_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _07526_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[0][26] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[1][26] ),
    .I2(\soc.spi_video_ram_1.write_fifo.fifo_mem[2][26] ),
    .I3(\soc.spi_video_ram_1.write_fifo.fifo_mem[3][26] ),
    .S0(_02919_),
    .S1(_02577_),
    .Z(_03174_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07527_ (.I(\soc.spi_video_ram_1.write_fifo.fifo_mem[7][26] ),
    .ZN(_03175_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07528_ (.A1(_02574_),
    .A2(_03175_),
    .ZN(_03176_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07529_ (.A1(_02700_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[6][26] ),
    .B(_03176_),
    .C(_02577_),
    .ZN(_03177_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07530_ (.I(\soc.spi_video_ram_1.write_fifo.fifo_mem[5][26] ),
    .ZN(_03178_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07531_ (.A1(_02919_),
    .A2(_03178_),
    .ZN(_03179_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07532_ (.A1(_02700_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[4][26] ),
    .B(_03179_),
    .C(_02741_),
    .ZN(_03180_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07533_ (.A1(_02706_),
    .A2(_03177_),
    .A3(_03180_),
    .ZN(_03181_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07534_ (.A1(_02984_),
    .A2(_03174_),
    .B(_03181_),
    .C(_02601_),
    .ZN(_03182_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07535_ (.A1(_03173_),
    .A2(_03182_),
    .B(_02567_),
    .ZN(_03183_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _07536_ (.A1(_02620_),
    .A2(_03165_),
    .B(_03183_),
    .C(_03019_),
    .ZN(_03184_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07537_ (.A1(_03146_),
    .A2(_03184_),
    .ZN(_03185_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07538_ (.A1(_01419_),
    .A2(_03107_),
    .B1(_03185_),
    .B2(_02677_),
    .ZN(_03186_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07539_ (.A1(\soc.spi_video_ram_1.output_buffer[11] ),
    .A2(_02676_),
    .ZN(_03187_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07540_ (.A1(_03015_),
    .A2(_03186_),
    .B(_03187_),
    .ZN(_00245_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07541_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[22][13] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[23][13] ),
    .S(_02700_),
    .Z(_03188_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07542_ (.I(\soc.spi_video_ram_1.write_fifo.fifo_mem[21][13] ),
    .ZN(_03189_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07543_ (.A1(_02591_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[20][13] ),
    .ZN(_03190_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _07544_ (.A1(_02764_),
    .A2(_03189_),
    .B(_03190_),
    .C(_02578_),
    .ZN(_03191_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _07545_ (.A1(_03041_),
    .A2(_03188_),
    .B(_03191_),
    .C(_02570_),
    .ZN(_03192_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07546_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[18][13] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[19][13] ),
    .S(_02651_),
    .Z(_03193_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07547_ (.A1(_02920_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[17][13] ),
    .ZN(_03194_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07548_ (.A1(_02926_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[16][13] ),
    .ZN(_03195_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07549_ (.A1(_03194_),
    .A2(_03195_),
    .B(_02976_),
    .ZN(_03196_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _07550_ (.A1(_02693_),
    .A2(_03193_),
    .B(_03196_),
    .C(_02984_),
    .ZN(_03197_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _07551_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[24][13] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[25][13] ),
    .I2(\soc.spi_video_ram_1.write_fifo.fifo_mem[26][13] ),
    .I3(\soc.spi_video_ram_1.write_fifo.fifo_mem[27][13] ),
    .S0(_03139_),
    .S1(_02908_),
    .Z(_03198_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07552_ (.I(\soc.spi_video_ram_1.write_fifo.fifo_mem[31][13] ),
    .ZN(_03199_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07553_ (.A1(_02907_),
    .A2(_03199_),
    .ZN(_03200_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07554_ (.A1(_02924_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[30][13] ),
    .B(_03200_),
    .C(_02908_),
    .ZN(_03201_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07555_ (.I(\soc.spi_video_ram_1.write_fifo.fifo_mem[29][13] ),
    .ZN(_03202_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07556_ (.A1(_02907_),
    .A2(_03202_),
    .ZN(_03203_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07557_ (.A1(_02924_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[28][13] ),
    .B(_03203_),
    .C(_02927_),
    .ZN(_03204_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07558_ (.A1(_02588_),
    .A2(_03201_),
    .A3(_03204_),
    .ZN(_03205_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07559_ (.A1(_02707_),
    .A2(_03198_),
    .B(_03205_),
    .C(_02970_),
    .ZN(_03206_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _07560_ (.A1(_02586_),
    .A2(_03192_),
    .A3(_03197_),
    .B(_03206_),
    .ZN(_03207_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07561_ (.A1(_02920_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[10][13] ),
    .ZN(_03208_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07562_ (.A1(_02922_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[11][13] ),
    .B(_02647_),
    .ZN(_03209_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07563_ (.I(\soc.spi_video_ram_1.write_fifo.fifo_mem[9][13] ),
    .ZN(_03210_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07564_ (.A1(_03139_),
    .A2(_03210_),
    .ZN(_03211_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07565_ (.A1(_02744_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[8][13] ),
    .B(_03211_),
    .ZN(_03212_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _07566_ (.A1(_03208_),
    .A2(_03209_),
    .B1(_03212_),
    .B2(_02976_),
    .C(_02929_),
    .ZN(_03213_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07567_ (.I(\soc.spi_video_ram_1.write_fifo.fifo_mem[15][13] ),
    .ZN(_03214_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07568_ (.A1(_02712_),
    .A2(_03214_),
    .ZN(_03215_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07569_ (.A1(_02784_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[14][13] ),
    .B(_03215_),
    .C(_02647_),
    .ZN(_03216_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _07570_ (.A1(_02919_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[12][13] ),
    .Z(_03217_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07571_ (.A1(_03021_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[13][13] ),
    .B(_03217_),
    .C(_03024_),
    .ZN(_03218_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07572_ (.A1(_02582_),
    .A2(_03216_),
    .A3(_03218_),
    .ZN(_03219_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07573_ (.A1(_02831_),
    .A2(_03213_),
    .A3(_03219_),
    .ZN(_03220_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _07574_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[0][13] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[1][13] ),
    .I2(\soc.spi_video_ram_1.write_fifo.fifo_mem[2][13] ),
    .I3(\soc.spi_video_ram_1.write_fifo.fifo_mem[3][13] ),
    .S0(_03139_),
    .S1(_02895_),
    .Z(_03221_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07575_ (.I(\soc.spi_video_ram_1.write_fifo.fifo_mem[7][13] ),
    .ZN(_03222_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07576_ (.A1(_02907_),
    .A2(_03222_),
    .ZN(_03223_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07577_ (.A1(_02924_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[6][13] ),
    .B(_03223_),
    .C(_02895_),
    .ZN(_03224_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07578_ (.I(\soc.spi_video_ram_1.write_fifo.fifo_mem[5][13] ),
    .ZN(_03225_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07579_ (.A1(_03139_),
    .A2(_03225_),
    .ZN(_03226_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07580_ (.A1(_02924_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[4][13] ),
    .B(_03226_),
    .C(_02927_),
    .ZN(_03227_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07581_ (.A1(_02582_),
    .A2(_03224_),
    .A3(_03227_),
    .ZN(_03228_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07582_ (.A1(_02707_),
    .A2(_03221_),
    .B(_03228_),
    .C(_02910_),
    .ZN(_03229_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07583_ (.A1(_02656_),
    .A2(_03220_),
    .A3(_03229_),
    .ZN(_03230_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07584_ (.A1(_02710_),
    .A2(_03207_),
    .B(_03230_),
    .C(_03019_),
    .ZN(_03231_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07585_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[18][25] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[19][25] ),
    .S(_02591_),
    .Z(_03232_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07586_ (.A1(_02920_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[17][25] ),
    .ZN(_03233_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07587_ (.A1(_02926_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[16][25] ),
    .ZN(_03234_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07588_ (.A1(_03233_),
    .A2(_03234_),
    .B(_02976_),
    .ZN(_03235_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _07589_ (.A1(_02693_),
    .A2(_03232_),
    .B(_03235_),
    .C(_02901_),
    .ZN(_03236_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07590_ (.I(\soc.spi_video_ram_1.write_fifo.fifo_mem[23][25] ),
    .ZN(_03237_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07591_ (.A1(_02591_),
    .A2(_03237_),
    .ZN(_03238_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07592_ (.A1(_02689_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[22][25] ),
    .B(_03238_),
    .C(_02598_),
    .ZN(_03239_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07593_ (.I(\soc.spi_video_ram_1.write_fifo.fifo_mem[21][25] ),
    .ZN(_03240_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07594_ (.A1(_02591_),
    .A2(_03240_),
    .ZN(_03241_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07595_ (.A1(_02689_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[20][25] ),
    .B(_03241_),
    .C(_02742_),
    .ZN(_03242_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07596_ (.A1(_02984_),
    .A2(_03239_),
    .A3(_03242_),
    .ZN(_03243_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07597_ (.A1(_02618_),
    .A2(_03243_),
    .ZN(_03244_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _07598_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[24][25] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[25][25] ),
    .I2(\soc.spi_video_ram_1.write_fifo.fifo_mem[26][25] ),
    .I3(\soc.spi_video_ram_1.write_fifo.fifo_mem[27][25] ),
    .S0(_02907_),
    .S1(_02908_),
    .Z(_03245_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07599_ (.I(\soc.spi_video_ram_1.write_fifo.fifo_mem[31][25] ),
    .ZN(_03246_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07600_ (.A1(_03054_),
    .A2(_03246_),
    .ZN(_03247_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07601_ (.A1(_02575_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[30][25] ),
    .B(_03247_),
    .C(_02904_),
    .ZN(_03248_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07602_ (.I(\soc.spi_video_ram_1.write_fifo.fifo_mem[29][25] ),
    .ZN(_03249_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07603_ (.A1(_03054_),
    .A2(_03249_),
    .ZN(_03250_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07604_ (.A1(_02575_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[28][25] ),
    .B(_03250_),
    .C(_02943_),
    .ZN(_03251_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07605_ (.A1(_02588_),
    .A2(_03248_),
    .A3(_03251_),
    .ZN(_03252_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07606_ (.A1(_02901_),
    .A2(_03245_),
    .B(_03252_),
    .C(_02970_),
    .ZN(_03253_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07607_ (.A1(_03236_),
    .A2(_03244_),
    .B(_03253_),
    .C(_02567_),
    .ZN(_03254_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _07608_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[0][25] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[1][25] ),
    .I2(\soc.spi_video_ram_1.write_fifo.fifo_mem[2][25] ),
    .I3(\soc.spi_video_ram_1.write_fifo.fifo_mem[3][25] ),
    .S0(_02680_),
    .S1(_02838_),
    .Z(_03255_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07609_ (.I(\soc.spi_video_ram_1.write_fifo.fifo_mem[5][25] ),
    .ZN(_03256_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07610_ (.A1(_02688_),
    .A2(_03256_),
    .ZN(_03257_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07611_ (.A1(_02920_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[4][25] ),
    .B(_03257_),
    .C(_03024_),
    .ZN(_03258_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07612_ (.I(\soc.spi_video_ram_1.write_fifo.fifo_mem[7][25] ),
    .ZN(_03259_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07613_ (.A1(_02763_),
    .A2(_03259_),
    .ZN(_03260_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07614_ (.A1(_02971_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[6][25] ),
    .B(_03260_),
    .C(_02838_),
    .ZN(_03261_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07615_ (.A1(_02582_),
    .A2(_03258_),
    .A3(_03261_),
    .ZN(_03262_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07616_ (.A1(_02767_),
    .A2(_03255_),
    .B(_03262_),
    .C(_02719_),
    .ZN(_03263_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07617_ (.A1(_03047_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[10][25] ),
    .ZN(_03264_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07618_ (.A1(_02704_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[11][25] ),
    .B(_02593_),
    .ZN(_03265_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07619_ (.I(\soc.spi_video_ram_1.write_fifo.fifo_mem[9][25] ),
    .ZN(_03266_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07620_ (.A1(_02763_),
    .A2(_03266_),
    .ZN(_03267_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07621_ (.A1(_02752_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[8][25] ),
    .B(_03267_),
    .ZN(_03268_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _07622_ (.A1(_03264_),
    .A2(_03265_),
    .B1(_03268_),
    .B2(_02691_),
    .C(_02929_),
    .ZN(_03269_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07623_ (.I(\soc.spi_video_ram_1.write_fifo.fifo_mem[15][25] ),
    .ZN(_03270_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07624_ (.A1(_02613_),
    .A2(_03270_),
    .ZN(_03271_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07625_ (.A1(_03047_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[14][25] ),
    .B(_03271_),
    .C(_02593_),
    .ZN(_03272_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _07626_ (.A1(_02931_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[12][25] ),
    .Z(_03273_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07627_ (.A1(_02704_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[13][25] ),
    .B(_03273_),
    .C(_02742_),
    .ZN(_03274_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07628_ (.A1(_02952_),
    .A2(_03272_),
    .A3(_03274_),
    .ZN(_03275_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07629_ (.A1(_02640_),
    .A2(_03269_),
    .A3(_03275_),
    .ZN(_03276_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07630_ (.A1(_02656_),
    .A2(_03263_),
    .A3(_03276_),
    .ZN(_03277_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07631_ (.A1(_02918_),
    .A2(_03254_),
    .A3(_03277_),
    .ZN(_03278_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07632_ (.A1(\soc.spi_video_ram_1.current_state[1] ),
    .A2(_02624_),
    .ZN(_03279_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07633_ (.A1(_03231_),
    .A2(_03278_),
    .B(_03279_),
    .ZN(_03280_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _07634_ (.A1(_02034_),
    .A2(_01897_),
    .A3(_02625_),
    .B(_02734_),
    .ZN(_03281_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _07635_ (.A1(\soc.spi_video_ram_1.output_buffer[10] ),
    .A2(_02882_),
    .B1(_03280_),
    .B2(_03281_),
    .ZN(_03282_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07636_ (.I(_03282_),
    .ZN(_00246_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07637_ (.A1(\soc.video_generator_1.v_count[3] ),
    .A2(_01897_),
    .ZN(_03283_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07638_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[18][14] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[19][14] ),
    .S(_02612_),
    .Z(_03284_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07639_ (.A1(_02931_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[17][14] ),
    .ZN(_03285_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07640_ (.A1(_02695_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[16][14] ),
    .ZN(_03286_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07641_ (.A1(_03285_),
    .A2(_03286_),
    .B(_02690_),
    .ZN(_03287_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _07642_ (.A1(_02958_),
    .A2(_03284_),
    .B(_03287_),
    .C(_02706_),
    .ZN(_03288_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07643_ (.A1(_02893_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[22][14] ),
    .ZN(_03289_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07644_ (.A1(_02703_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[23][14] ),
    .B(_02592_),
    .ZN(_03290_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07645_ (.I(\soc.spi_video_ram_1.write_fifo.fifo_mem[21][14] ),
    .ZN(_03291_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07646_ (.A1(_02679_),
    .A2(_03291_),
    .ZN(_03292_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07647_ (.A1(_02783_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[20][14] ),
    .B(_03292_),
    .C(_02741_),
    .ZN(_03293_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07648_ (.A1(_03289_),
    .A2(_03290_),
    .B(_03293_),
    .C(_02581_),
    .ZN(_03294_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07649_ (.A1(_02601_),
    .A2(_03294_),
    .ZN(_03295_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _07650_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[24][14] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[25][14] ),
    .I2(\soc.spi_video_ram_1.write_fifo.fifo_mem[26][14] ),
    .I3(\soc.spi_video_ram_1.write_fifo.fifo_mem[27][14] ),
    .S0(_02902_),
    .S1(_02894_),
    .Z(_03296_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07651_ (.I(\soc.spi_video_ram_1.write_fifo.fifo_mem[31][14] ),
    .ZN(_03297_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07652_ (.A1(_02902_),
    .A2(_03297_),
    .ZN(_03298_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07653_ (.A1(_02574_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[30][14] ),
    .B(_03298_),
    .C(_02894_),
    .ZN(_03299_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07654_ (.I(\soc.spi_video_ram_1.write_fifo.fifo_mem[29][14] ),
    .ZN(_03300_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07655_ (.A1(_02902_),
    .A2(_03300_),
    .ZN(_03301_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07656_ (.A1(_02574_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[28][14] ),
    .B(_03301_),
    .C(_02741_),
    .ZN(_03302_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07657_ (.A1(_02581_),
    .A2(_03299_),
    .A3(_03302_),
    .ZN(_03303_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07658_ (.A1(_02642_),
    .A2(_03296_),
    .B(_03303_),
    .C(_02585_),
    .ZN(_03304_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07659_ (.A1(_03288_),
    .A2(_03295_),
    .B(_03304_),
    .ZN(_03305_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07660_ (.A1(_02783_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[10][14] ),
    .ZN(_03306_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07661_ (.A1(_02695_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[11][14] ),
    .B(_02894_),
    .ZN(_03307_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07662_ (.I(\soc.spi_video_ram_1.write_fifo.fifo_mem[9][14] ),
    .ZN(_03308_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07663_ (.A1(_02902_),
    .A2(_03308_),
    .ZN(_03309_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07664_ (.A1(_02590_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[8][14] ),
    .B(_03309_),
    .ZN(_03310_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _07665_ (.A1(_03306_),
    .A2(_03307_),
    .B1(_03310_),
    .B2(_02690_),
    .C(_02569_),
    .ZN(_03311_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07666_ (.I(\soc.spi_video_ram_1.write_fifo.fifo_mem[15][14] ),
    .ZN(_03312_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07667_ (.A1(_02644_),
    .A2(_03312_),
    .ZN(_03313_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07668_ (.A1(_02931_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[14][14] ),
    .B(_03313_),
    .C(_02646_),
    .ZN(_03314_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _07669_ (.A1(_02573_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[12][14] ),
    .Z(_03315_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07670_ (.A1(_02695_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[13][14] ),
    .B(_03315_),
    .C(_02741_),
    .ZN(_03316_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07671_ (.A1(_02581_),
    .A2(_03314_),
    .A3(_03316_),
    .ZN(_03317_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07672_ (.A1(_02585_),
    .A2(_03311_),
    .A3(_03317_),
    .ZN(_03318_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _07673_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[0][14] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[1][14] ),
    .I2(\soc.spi_video_ram_1.write_fifo.fifo_mem[2][14] ),
    .I3(\soc.spi_video_ram_1.write_fifo.fifo_mem[3][14] ),
    .S0(_02902_),
    .S1(_02894_),
    .Z(_03319_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07674_ (.I(\soc.spi_video_ram_1.write_fifo.fifo_mem[5][14] ),
    .ZN(_03320_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07675_ (.A1(_02902_),
    .A2(_03320_),
    .ZN(_03321_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07676_ (.A1(_02574_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[4][14] ),
    .B(_03321_),
    .C(_02740_),
    .ZN(_03322_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07677_ (.I(\soc.spi_video_ram_1.write_fifo.fifo_mem[7][14] ),
    .ZN(_03323_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07678_ (.A1(_02902_),
    .A2(_03323_),
    .ZN(_03324_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07679_ (.A1(_02574_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[6][14] ),
    .B(_03324_),
    .C(_02894_),
    .ZN(_03325_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07680_ (.A1(_02581_),
    .A2(_03322_),
    .A3(_03325_),
    .ZN(_03326_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07681_ (.A1(_02706_),
    .A2(_03319_),
    .B(_03326_),
    .C(_02600_),
    .ZN(_03327_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07682_ (.A1(_02655_),
    .A2(_03318_),
    .A3(_03327_),
    .ZN(_03328_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07683_ (.A1(_02655_),
    .A2(_03305_),
    .B(_03328_),
    .ZN(_03329_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07684_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[18][24] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[19][24] ),
    .S(_02612_),
    .Z(_03330_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07685_ (.A1(_02783_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[17][24] ),
    .ZN(_03331_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07686_ (.A1(_02695_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[16][24] ),
    .ZN(_03332_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07687_ (.A1(_03331_),
    .A2(_03332_),
    .B(_02577_),
    .ZN(_03333_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _07688_ (.A1(_02958_),
    .A2(_03330_),
    .B(_03333_),
    .C(_02706_),
    .ZN(_03334_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07689_ (.I(\soc.spi_video_ram_1.write_fifo.fifo_mem[23][24] ),
    .ZN(_03335_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07690_ (.A1(_02612_),
    .A2(_03335_),
    .ZN(_03336_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07691_ (.A1(_02893_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[22][24] ),
    .B(_03336_),
    .C(_02592_),
    .ZN(_03337_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07692_ (.I(\soc.spi_video_ram_1.write_fifo.fifo_mem[21][24] ),
    .ZN(_03338_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07693_ (.A1(_02612_),
    .A2(_03338_),
    .ZN(_03339_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07694_ (.A1(_02893_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[20][24] ),
    .B(_03339_),
    .C(_02741_),
    .ZN(_03340_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07695_ (.A1(_02900_),
    .A2(_03337_),
    .A3(_03340_),
    .ZN(_03341_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07696_ (.A1(_02601_),
    .A2(_03341_),
    .ZN(_03342_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _07697_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[24][24] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[25][24] ),
    .I2(\soc.spi_video_ram_1.write_fifo.fifo_mem[26][24] ),
    .I3(\soc.spi_video_ram_1.write_fifo.fifo_mem[27][24] ),
    .S0(_02902_),
    .S1(_02576_),
    .Z(_03343_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07698_ (.I(\soc.spi_video_ram_1.write_fifo.fifo_mem[31][24] ),
    .ZN(_03344_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07699_ (.A1(_02573_),
    .A2(_03344_),
    .ZN(_03345_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07700_ (.A1(_02590_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[30][24] ),
    .B(_03345_),
    .C(_02576_),
    .ZN(_03346_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07701_ (.I(\soc.spi_video_ram_1.write_fifo.fifo_mem[29][24] ),
    .ZN(_03347_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07702_ (.A1(_02573_),
    .A2(_03347_),
    .ZN(_03348_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07703_ (.A1(_02590_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[28][24] ),
    .B(_03348_),
    .C(_02740_),
    .ZN(_03349_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07704_ (.A1(_02581_),
    .A2(_03346_),
    .A3(_03349_),
    .ZN(_03350_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07705_ (.A1(_02706_),
    .A2(_03343_),
    .B(_03350_),
    .C(_00003_),
    .ZN(_03351_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07706_ (.A1(_03334_),
    .A2(_03342_),
    .B(_03351_),
    .C(_00004_),
    .ZN(_03352_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _07707_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[0][24] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[1][24] ),
    .I2(\soc.spi_video_ram_1.write_fifo.fifo_mem[2][24] ),
    .I3(\soc.spi_video_ram_1.write_fifo.fifo_mem[3][24] ),
    .S0(_02679_),
    .S1(_02894_),
    .Z(_03353_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07708_ (.I(\soc.spi_video_ram_1.write_fifo.fifo_mem[7][24] ),
    .ZN(_03354_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07709_ (.A1(_02679_),
    .A2(_03354_),
    .ZN(_03355_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07710_ (.A1(_02783_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[6][24] ),
    .B(_03355_),
    .C(_02894_),
    .ZN(_03356_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07711_ (.I(\soc.spi_video_ram_1.write_fifo.fifo_mem[5][24] ),
    .ZN(_03357_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07712_ (.A1(_02679_),
    .A2(_03357_),
    .ZN(_03358_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07713_ (.A1(_02783_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[4][24] ),
    .B(_03358_),
    .C(_02741_),
    .ZN(_03359_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07714_ (.A1(_02581_),
    .A2(_03356_),
    .A3(_03359_),
    .ZN(_03360_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07715_ (.A1(_02642_),
    .A2(_03353_),
    .B(_03360_),
    .C(_02601_),
    .ZN(_03361_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07716_ (.A1(_02903_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[10][24] ),
    .ZN(_03362_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07717_ (.A1(_02703_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[11][24] ),
    .B(_02646_),
    .ZN(_03363_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07718_ (.I(\soc.spi_video_ram_1.write_fifo.fifo_mem[9][24] ),
    .ZN(_03364_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07719_ (.A1(_02679_),
    .A2(_03364_),
    .ZN(_03365_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07720_ (.A1(_02919_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[8][24] ),
    .B(_03365_),
    .ZN(_03366_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _07721_ (.A1(_03362_),
    .A2(_03363_),
    .B1(_03366_),
    .B2(_02908_),
    .C(_02569_),
    .ZN(_03367_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07722_ (.I(\soc.spi_video_ram_1.write_fifo.fifo_mem[15][24] ),
    .ZN(_03368_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07723_ (.A1(_02644_),
    .A2(_03368_),
    .ZN(_03369_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07724_ (.A1(_03139_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[14][24] ),
    .B(_03369_),
    .C(_02646_),
    .ZN(_03370_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _07725_ (.A1(_02573_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[12][24] ),
    .Z(_03371_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07726_ (.A1(_02703_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[13][24] ),
    .B(_03371_),
    .C(_02741_),
    .ZN(_03372_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07727_ (.A1(_02900_),
    .A2(_03370_),
    .A3(_03372_),
    .ZN(_03373_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07728_ (.A1(_02585_),
    .A2(_03367_),
    .A3(_03373_),
    .ZN(_03374_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07729_ (.A1(_02655_),
    .A2(_03361_),
    .A3(_03374_),
    .ZN(_03375_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07730_ (.A1(_03352_),
    .A2(_03375_),
    .ZN(_03376_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07731_ (.I0(_03329_),
    .I1(_03376_),
    .S(_02918_),
    .Z(_03377_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _07732_ (.A1(_03283_),
    .A2(_02625_),
    .B1(_03279_),
    .B2(_03377_),
    .C(_02734_),
    .ZN(_03378_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07733_ (.A1(\soc.spi_video_ram_1.output_buffer[9] ),
    .A2(_02882_),
    .B(_03378_),
    .ZN(_03379_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07734_ (.I(_03379_),
    .ZN(_00247_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07735_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[18][15] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[19][15] ),
    .S(_02597_),
    .Z(_03380_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07736_ (.A1(_03047_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[17][15] ),
    .ZN(_03381_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07737_ (.A1(_02922_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[16][15] ),
    .ZN(_03382_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07738_ (.A1(_03381_),
    .A2(_03382_),
    .B(_02976_),
    .ZN(_03383_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _07739_ (.A1(_02693_),
    .A2(_03380_),
    .B(_03383_),
    .C(_02707_),
    .ZN(_03384_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07740_ (.A1(_02764_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[22][15] ),
    .ZN(_03385_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07741_ (.A1(_02704_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[23][15] ),
    .B(_02958_),
    .ZN(_03386_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07742_ (.I(\soc.spi_video_ram_1.write_fifo.fifo_mem[21][15] ),
    .ZN(_03387_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07743_ (.A1(_02712_),
    .A2(_03387_),
    .ZN(_03388_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07744_ (.A1(_02784_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[20][15] ),
    .B(_03388_),
    .C(_03024_),
    .ZN(_03389_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07745_ (.A1(_03385_),
    .A2(_03386_),
    .B(_03389_),
    .C(_02952_),
    .ZN(_03390_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07746_ (.A1(_02602_),
    .A2(_03390_),
    .ZN(_03391_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _07747_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[24][15] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[25][15] ),
    .I2(\soc.spi_video_ram_1.write_fifo.fifo_mem[26][15] ),
    .I3(\soc.spi_video_ram_1.write_fifo.fifo_mem[27][15] ),
    .S0(_02688_),
    .S1(_02827_),
    .Z(_03392_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07748_ (.I(\soc.spi_video_ram_1.write_fifo.fifo_mem[31][15] ),
    .ZN(_03393_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07749_ (.A1(_02893_),
    .A2(_03393_),
    .ZN(_03394_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07750_ (.A1(_02752_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[30][15] ),
    .B(_03394_),
    .C(_02827_),
    .ZN(_03395_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07751_ (.I(\soc.spi_video_ram_1.write_fifo.fifo_mem[29][15] ),
    .ZN(_03396_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07752_ (.A1(_02893_),
    .A2(_03396_),
    .ZN(_03397_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07753_ (.A1(_02752_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[28][15] ),
    .B(_03397_),
    .C(_02927_),
    .ZN(_03398_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07754_ (.A1(_02582_),
    .A2(_03395_),
    .A3(_03398_),
    .ZN(_03399_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07755_ (.A1(_02767_),
    .A2(_03392_),
    .B(_03399_),
    .C(_02970_),
    .ZN(_03400_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07756_ (.A1(_03384_),
    .A2(_03391_),
    .B(_03400_),
    .ZN(_03401_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _07757_ (.A1(_02919_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[12][15] ),
    .Z(_03402_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07758_ (.A1(_03021_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[13][15] ),
    .B(_03402_),
    .C(_03024_),
    .ZN(_03403_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07759_ (.I(\soc.spi_video_ram_1.write_fifo.fifo_mem[15][15] ),
    .ZN(_03404_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07760_ (.A1(_02712_),
    .A2(_03404_),
    .ZN(_03405_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07761_ (.A1(_02784_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[14][15] ),
    .B(_03405_),
    .C(_02647_),
    .ZN(_03406_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07762_ (.A1(_02952_),
    .A2(_03403_),
    .A3(_03406_),
    .ZN(_03407_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07763_ (.A1(_02920_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[10][15] ),
    .ZN(_03408_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07764_ (.A1(_02922_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[11][15] ),
    .B(_02647_),
    .ZN(_03409_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07765_ (.I(\soc.spi_video_ram_1.write_fifo.fifo_mem[9][15] ),
    .ZN(_03410_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07766_ (.A1(_03139_),
    .A2(_03410_),
    .ZN(_03411_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07767_ (.A1(_02744_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[8][15] ),
    .B(_03411_),
    .ZN(_03412_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _07768_ (.A1(_03408_),
    .A2(_03409_),
    .B1(_03412_),
    .B2(_02976_),
    .C(_02929_),
    .ZN(_03413_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07769_ (.A1(_02831_),
    .A2(_03407_),
    .A3(_03413_),
    .ZN(_03414_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _07770_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[0][15] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[1][15] ),
    .I2(\soc.spi_video_ram_1.write_fifo.fifo_mem[2][15] ),
    .I3(\soc.spi_video_ram_1.write_fifo.fifo_mem[3][15] ),
    .S0(_03139_),
    .S1(_02895_),
    .Z(_03415_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07771_ (.I(\soc.spi_video_ram_1.write_fifo.fifo_mem[7][15] ),
    .ZN(_03416_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07772_ (.A1(_02907_),
    .A2(_03416_),
    .ZN(_03417_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07773_ (.A1(_02924_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[6][15] ),
    .B(_03417_),
    .C(_02895_),
    .ZN(_03418_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07774_ (.I(\soc.spi_video_ram_1.write_fifo.fifo_mem[5][15] ),
    .ZN(_03419_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07775_ (.A1(_02907_),
    .A2(_03419_),
    .ZN(_03420_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07776_ (.A1(_02924_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[4][15] ),
    .B(_03420_),
    .C(_02927_),
    .ZN(_03421_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07777_ (.A1(_02588_),
    .A2(_03418_),
    .A3(_03421_),
    .ZN(_03422_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07778_ (.A1(_02707_),
    .A2(_03415_),
    .B(_03422_),
    .C(_02910_),
    .ZN(_03423_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07779_ (.A1(_02656_),
    .A2(_03414_),
    .A3(_03423_),
    .ZN(_03424_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07780_ (.A1(_02656_),
    .A2(_03401_),
    .B(_03424_),
    .C(_03019_),
    .ZN(_03425_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07781_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[18][23] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[19][23] ),
    .S(_02591_),
    .Z(_03426_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07782_ (.A1(_02920_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[17][23] ),
    .ZN(_03427_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07783_ (.A1(_02926_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[16][23] ),
    .ZN(_03428_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07784_ (.A1(_03427_),
    .A2(_03428_),
    .B(_02976_),
    .ZN(_03429_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _07785_ (.A1(_02693_),
    .A2(_03426_),
    .B(_03429_),
    .C(_02901_),
    .ZN(_03430_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07786_ (.I(\soc.spi_video_ram_1.write_fifo.fifo_mem[23][23] ),
    .ZN(_03431_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07787_ (.A1(_02591_),
    .A2(_03431_),
    .ZN(_03432_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07788_ (.A1(_02689_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[22][23] ),
    .B(_03432_),
    .C(_02598_),
    .ZN(_03433_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07789_ (.I(\soc.spi_video_ram_1.write_fifo.fifo_mem[21][23] ),
    .ZN(_03434_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07790_ (.A1(_02651_),
    .A2(_03434_),
    .ZN(_03435_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07791_ (.A1(_02689_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[20][23] ),
    .B(_03435_),
    .C(_02742_),
    .ZN(_03436_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07792_ (.A1(_02984_),
    .A2(_03433_),
    .A3(_03436_),
    .ZN(_03437_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07793_ (.A1(_02618_),
    .A2(_03437_),
    .ZN(_03438_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _07794_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[24][23] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[25][23] ),
    .I2(\soc.spi_video_ram_1.write_fifo.fifo_mem[26][23] ),
    .I3(\soc.spi_video_ram_1.write_fifo.fifo_mem[27][23] ),
    .S0(_02903_),
    .S1(_02904_),
    .Z(_03439_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07795_ (.I(\soc.spi_video_ram_1.write_fifo.fifo_mem[31][23] ),
    .ZN(_03440_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07796_ (.A1(_03054_),
    .A2(_03440_),
    .ZN(_03441_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07797_ (.A1(_02575_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[30][23] ),
    .B(_03441_),
    .C(_02904_),
    .ZN(_03442_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07798_ (.I(\soc.spi_video_ram_1.write_fifo.fifo_mem[29][23] ),
    .ZN(_03443_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07799_ (.A1(_03054_),
    .A2(_03443_),
    .ZN(_03444_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07800_ (.A1(_02575_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[28][23] ),
    .B(_03444_),
    .C(_02943_),
    .ZN(_03445_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07801_ (.A1(_02588_),
    .A2(_03442_),
    .A3(_03445_),
    .ZN(_03446_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07802_ (.A1(_02901_),
    .A2(_03439_),
    .B(_03446_),
    .C(_02970_),
    .ZN(_03447_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07803_ (.A1(_03430_),
    .A2(_03438_),
    .B(_03447_),
    .C(_02567_),
    .ZN(_03448_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _07804_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[0][23] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[1][23] ),
    .I2(\soc.spi_video_ram_1.write_fifo.fifo_mem[2][23] ),
    .I3(\soc.spi_video_ram_1.write_fifo.fifo_mem[3][23] ),
    .S0(_02680_),
    .S1(_02838_),
    .Z(_03449_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07805_ (.I(\soc.spi_video_ram_1.write_fifo.fifo_mem[7][23] ),
    .ZN(_03450_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07806_ (.A1(_02688_),
    .A2(_03450_),
    .ZN(_03451_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07807_ (.A1(_02920_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[6][23] ),
    .B(_03451_),
    .C(_02838_),
    .ZN(_03452_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07808_ (.I(\soc.spi_video_ram_1.write_fifo.fifo_mem[5][23] ),
    .ZN(_03453_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07809_ (.A1(_02688_),
    .A2(_03453_),
    .ZN(_03454_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07810_ (.A1(_02971_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[4][23] ),
    .B(_03454_),
    .C(_03024_),
    .ZN(_03455_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07811_ (.A1(_02582_),
    .A2(_03452_),
    .A3(_03455_),
    .ZN(_03456_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07812_ (.A1(_02767_),
    .A2(_03449_),
    .B(_03456_),
    .C(_02719_),
    .ZN(_03457_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07813_ (.A1(_03047_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[10][23] ),
    .ZN(_03458_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07814_ (.A1(_02704_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[11][23] ),
    .B(_02593_),
    .ZN(_03459_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07815_ (.I(\soc.spi_video_ram_1.write_fifo.fifo_mem[9][23] ),
    .ZN(_03460_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07816_ (.A1(_02763_),
    .A2(_03460_),
    .ZN(_03461_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07817_ (.A1(_02752_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[8][23] ),
    .B(_03461_),
    .ZN(_03462_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _07818_ (.A1(_03458_),
    .A2(_03459_),
    .B1(_03462_),
    .B2(_02691_),
    .C(_02929_),
    .ZN(_03463_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07819_ (.I(\soc.spi_video_ram_1.write_fifo.fifo_mem[15][23] ),
    .ZN(_03464_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07820_ (.A1(_02613_),
    .A2(_03464_),
    .ZN(_03465_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07821_ (.A1(_03047_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[14][23] ),
    .B(_03465_),
    .C(_02593_),
    .ZN(_03466_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _07822_ (.A1(_02931_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[12][23] ),
    .Z(_03467_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07823_ (.A1(_02704_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[13][23] ),
    .B(_03467_),
    .C(_02742_),
    .ZN(_03468_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07824_ (.A1(_02952_),
    .A2(_03466_),
    .A3(_03468_),
    .ZN(_03469_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07825_ (.A1(_02640_),
    .A2(_03463_),
    .A3(_03469_),
    .ZN(_03470_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07826_ (.A1(_02656_),
    .A2(_03457_),
    .A3(_03470_),
    .ZN(_03471_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07827_ (.A1(_02918_),
    .A2(_03448_),
    .A3(_03471_),
    .ZN(_03472_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07828_ (.A1(_03425_),
    .A2(_03472_),
    .B(_03279_),
    .ZN(_03473_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07829_ (.A1(\soc.video_generator_1.v_count[2] ),
    .A2(_01897_),
    .ZN(_03474_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07830_ (.A1(_03474_),
    .A2(_02625_),
    .B(_02882_),
    .ZN(_03475_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _07831_ (.A1(\soc.spi_video_ram_1.output_buffer[8] ),
    .A2(_02882_),
    .B1(_03473_),
    .B2(_03475_),
    .ZN(_03476_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07832_ (.I(_03476_),
    .ZN(_00248_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07833_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[18][22] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[19][22] ),
    .S(_02575_),
    .Z(_03477_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07834_ (.A1(_03047_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[17][22] ),
    .ZN(_03478_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07835_ (.A1(_03021_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[16][22] ),
    .ZN(_03479_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07836_ (.A1(_03478_),
    .A2(_03479_),
    .B(_02976_),
    .ZN(_03480_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _07837_ (.A1(_02693_),
    .A2(_03477_),
    .B(_03480_),
    .C(_02707_),
    .ZN(_03481_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07838_ (.I(\soc.spi_video_ram_1.write_fifo.fifo_mem[23][22] ),
    .ZN(_03482_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07839_ (.A1(_02607_),
    .A2(_03482_),
    .ZN(_03483_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07840_ (.A1(_02764_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[22][22] ),
    .B(_03483_),
    .C(_02958_),
    .ZN(_03484_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07841_ (.I(\soc.spi_video_ram_1.write_fifo.fifo_mem[21][22] ),
    .ZN(_03485_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07842_ (.A1(_02607_),
    .A2(_03485_),
    .ZN(_03486_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07843_ (.A1(_02764_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[20][22] ),
    .B(_03486_),
    .C(_02742_),
    .ZN(_03487_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07844_ (.A1(_02984_),
    .A2(_03484_),
    .A3(_03487_),
    .ZN(_03488_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07845_ (.A1(_02602_),
    .A2(_03488_),
    .ZN(_03489_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _07846_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[24][22] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[25][22] ),
    .I2(\soc.spi_video_ram_1.write_fifo.fifo_mem[26][22] ),
    .I3(\soc.spi_video_ram_1.write_fifo.fifo_mem[27][22] ),
    .S0(_02893_),
    .S1(_02895_),
    .Z(_03490_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07847_ (.I(\soc.spi_video_ram_1.write_fifo.fifo_mem[31][22] ),
    .ZN(_03491_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07848_ (.A1(_03139_),
    .A2(_03491_),
    .ZN(_03492_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07849_ (.A1(_02752_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[30][22] ),
    .B(_03492_),
    .C(_02895_),
    .ZN(_03493_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07850_ (.I(\soc.spi_video_ram_1.write_fifo.fifo_mem[29][22] ),
    .ZN(_03494_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07851_ (.A1(_03139_),
    .A2(_03494_),
    .ZN(_03495_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07852_ (.A1(_02752_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[28][22] ),
    .B(_03495_),
    .C(_02927_),
    .ZN(_03496_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07853_ (.A1(_02582_),
    .A2(_03493_),
    .A3(_03496_),
    .ZN(_03497_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07854_ (.A1(_02767_),
    .A2(_03490_),
    .B(_03497_),
    .C(_02970_),
    .ZN(_03498_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07855_ (.A1(_03481_),
    .A2(_03489_),
    .B(_03498_),
    .C(_02567_),
    .ZN(_03499_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _07856_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[0][22] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[1][22] ),
    .I2(\soc.spi_video_ram_1.write_fifo.fifo_mem[2][22] ),
    .I3(\soc.spi_video_ram_1.write_fifo.fifo_mem[3][22] ),
    .S0(_02700_),
    .S1(_02647_),
    .Z(_03500_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07857_ (.I(\soc.spi_video_ram_1.write_fifo.fifo_mem[7][22] ),
    .ZN(_03501_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07858_ (.A1(_02700_),
    .A2(_03501_),
    .ZN(_03502_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07859_ (.A1(_03047_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[6][22] ),
    .B(_03502_),
    .C(_02647_),
    .ZN(_03503_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07860_ (.I(\soc.spi_video_ram_1.write_fifo.fifo_mem[5][22] ),
    .ZN(_03504_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07861_ (.A1(_02700_),
    .A2(_03504_),
    .ZN(_03505_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07862_ (.A1(_03047_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[4][22] ),
    .B(_03505_),
    .C(_03024_),
    .ZN(_03506_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07863_ (.A1(_02952_),
    .A2(_03503_),
    .A3(_03506_),
    .ZN(_03507_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07864_ (.A1(_02643_),
    .A2(_03500_),
    .B(_03507_),
    .C(_02719_),
    .ZN(_03508_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _07865_ (.A1(_02907_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[12][22] ),
    .Z(_03509_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07866_ (.A1(_02704_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[13][22] ),
    .B(_03509_),
    .C(_02742_),
    .ZN(_03510_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07867_ (.I(\soc.spi_video_ram_1.write_fifo.fifo_mem[15][22] ),
    .ZN(_03511_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07868_ (.A1(_02635_),
    .A2(_03511_),
    .ZN(_03512_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07869_ (.A1(_02764_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[14][22] ),
    .B(_03512_),
    .C(_02958_),
    .ZN(_03513_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07870_ (.A1(_02984_),
    .A2(_03510_),
    .A3(_03513_),
    .ZN(_03514_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07871_ (.A1(_02689_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[10][22] ),
    .ZN(_03515_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07872_ (.A1(_02704_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[11][22] ),
    .B(_02578_),
    .ZN(_03516_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07873_ (.I(\soc.spi_video_ram_1.write_fifo.fifo_mem[9][22] ),
    .ZN(_03517_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07874_ (.A1(_02712_),
    .A2(_03517_),
    .ZN(_03518_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07875_ (.A1(_02784_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[8][22] ),
    .B(_03518_),
    .ZN(_03519_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _07876_ (.A1(_03515_),
    .A2(_03516_),
    .B1(_03519_),
    .B2(_02723_),
    .C(_02570_),
    .ZN(_03520_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07877_ (.A1(_02640_),
    .A2(_03514_),
    .A3(_03520_),
    .ZN(_03521_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07878_ (.A1(_02656_),
    .A2(_03508_),
    .A3(_03521_),
    .ZN(_03522_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _07879_ (.A1(_02677_),
    .A2(_02918_),
    .A3(_03499_),
    .A4(_03522_),
    .ZN(_03523_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07880_ (.A1(_01885_),
    .A2(_02625_),
    .B(_03523_),
    .ZN(_03524_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07881_ (.I0(\soc.spi_video_ram_1.output_buffer[7] ),
    .I1(_03524_),
    .S(_02633_),
    .Z(_03525_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07882_ (.I(_03525_),
    .Z(_00249_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _07883_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[0][21] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[1][21] ),
    .I2(\soc.spi_video_ram_1.write_fifo.fifo_mem[2][21] ),
    .I3(\soc.spi_video_ram_1.write_fifo.fifo_mem[3][21] ),
    .S0(_02763_),
    .S1(_02827_),
    .Z(_03526_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07884_ (.I(\soc.spi_video_ram_1.write_fifo.fifo_mem[7][21] ),
    .ZN(_03527_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07885_ (.A1(_02688_),
    .A2(_03527_),
    .ZN(_03528_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07886_ (.A1(_02971_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[6][21] ),
    .B(_03528_),
    .C(_02827_),
    .ZN(_03529_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07887_ (.I(\soc.spi_video_ram_1.write_fifo.fifo_mem[5][21] ),
    .ZN(_03530_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07888_ (.A1(_02688_),
    .A2(_03530_),
    .ZN(_03531_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07889_ (.A1(_02971_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[4][21] ),
    .B(_03531_),
    .C(_02927_),
    .ZN(_03532_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07890_ (.A1(_02582_),
    .A2(_03529_),
    .A3(_03532_),
    .ZN(_03533_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07891_ (.A1(_02767_),
    .A2(_03526_),
    .B(_03533_),
    .C(_02910_),
    .ZN(_03534_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07892_ (.A1(_02784_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[10][21] ),
    .ZN(_03535_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07893_ (.A1(_03021_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[11][21] ),
    .B(_02652_),
    .ZN(_03536_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07894_ (.I(\soc.spi_video_ram_1.write_fifo.fifo_mem[9][21] ),
    .ZN(_03537_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07895_ (.A1(_02688_),
    .A2(_03537_),
    .ZN(_03538_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07896_ (.A1(_02752_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[8][21] ),
    .B(_03538_),
    .ZN(_03539_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _07897_ (.A1(_03535_),
    .A2(_03536_),
    .B1(_03539_),
    .B2(_02691_),
    .C(_02929_),
    .ZN(_03540_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07898_ (.I(\soc.spi_video_ram_1.write_fifo.fifo_mem[15][21] ),
    .ZN(_03541_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07899_ (.A1(_02645_),
    .A2(_03541_),
    .ZN(_03542_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07900_ (.A1(_03047_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[14][21] ),
    .B(_03542_),
    .C(_02652_),
    .ZN(_03543_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _07901_ (.A1(_02783_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[12][21] ),
    .Z(_03544_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07902_ (.A1(_02704_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[13][21] ),
    .B(_03544_),
    .C(_02742_),
    .ZN(_03545_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07903_ (.A1(_02952_),
    .A2(_03543_),
    .A3(_03545_),
    .ZN(_03546_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07904_ (.A1(_02831_),
    .A2(_03540_),
    .A3(_03546_),
    .ZN(_03547_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07905_ (.A1(_02656_),
    .A2(_03534_),
    .A3(_03547_),
    .ZN(_03548_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07906_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[18][21] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[19][21] ),
    .S(_02651_),
    .Z(_03549_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07907_ (.A1(_02920_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[17][21] ),
    .ZN(_03550_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07908_ (.A1(_02926_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[16][21] ),
    .ZN(_03551_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07909_ (.A1(_03550_),
    .A2(_03551_),
    .B(_02976_),
    .ZN(_03552_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _07910_ (.A1(_02693_),
    .A2(_03549_),
    .B(_03552_),
    .C(_02984_),
    .ZN(_03553_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07911_ (.I(\soc.spi_video_ram_1.write_fifo.fifo_mem[23][21] ),
    .ZN(_03554_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07912_ (.A1(_02651_),
    .A2(_03554_),
    .ZN(_03555_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07913_ (.A1(_02689_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[22][21] ),
    .B(_03555_),
    .C(_02593_),
    .ZN(_03556_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07914_ (.I(\soc.spi_video_ram_1.write_fifo.fifo_mem[21][21] ),
    .ZN(_03557_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07915_ (.A1(_02613_),
    .A2(_03557_),
    .ZN(_03558_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07916_ (.A1(_02689_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[20][21] ),
    .B(_03558_),
    .C(_02742_),
    .ZN(_03559_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07917_ (.A1(_02952_),
    .A2(_03556_),
    .A3(_03559_),
    .ZN(_03560_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07918_ (.A1(_02719_),
    .A2(_03560_),
    .ZN(_03561_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _07919_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[24][21] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[25][21] ),
    .I2(\soc.spi_video_ram_1.write_fifo.fifo_mem[26][21] ),
    .I3(\soc.spi_video_ram_1.write_fifo.fifo_mem[27][21] ),
    .S0(_02903_),
    .S1(_02904_),
    .Z(_03562_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07920_ (.I(\soc.spi_video_ram_1.write_fifo.fifo_mem[29][21] ),
    .ZN(_03563_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07921_ (.A1(_02931_),
    .A2(_03563_),
    .ZN(_03564_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07922_ (.A1(_02635_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[28][21] ),
    .B(_03564_),
    .C(_02943_),
    .ZN(_03565_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07923_ (.I(\soc.spi_video_ram_1.write_fifo.fifo_mem[31][21] ),
    .ZN(_03566_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07924_ (.A1(_02931_),
    .A2(_03566_),
    .ZN(_03567_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07925_ (.A1(_02635_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[30][21] ),
    .B(_03567_),
    .C(_02904_),
    .ZN(_03568_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07926_ (.A1(_02642_),
    .A2(_03565_),
    .A3(_03568_),
    .ZN(_03569_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07927_ (.A1(_02901_),
    .A2(_03562_),
    .B(_03569_),
    .C(_02970_),
    .ZN(_03570_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07928_ (.A1(_03553_),
    .A2(_03561_),
    .B(_03570_),
    .C(_02567_),
    .ZN(_03571_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _07929_ (.A1(_02677_),
    .A2(_01392_),
    .A3(_03548_),
    .A4(_03571_),
    .ZN(_03572_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07930_ (.A1(_01898_),
    .A2(_02625_),
    .B(_03572_),
    .C(_02734_),
    .ZN(_03573_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07931_ (.A1(\soc.spi_video_ram_1.output_buffer[6] ),
    .A2(_02882_),
    .B(_03573_),
    .ZN(_03574_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07932_ (.I(_03574_),
    .ZN(_00250_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _07933_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[8][20] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[9][20] ),
    .I2(\soc.spi_video_ram_1.write_fifo.fifo_mem[10][20] ),
    .I3(\soc.spi_video_ram_1.write_fifo.fifo_mem[11][20] ),
    .S0(_02717_),
    .S1(_02682_),
    .Z(_03575_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07934_ (.A1(_02678_),
    .A2(_03575_),
    .ZN(_03576_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07935_ (.I(_02596_),
    .Z(_03577_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _07936_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[12][20] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[13][20] ),
    .I2(\soc.spi_video_ram_1.write_fifo.fifo_mem[14][20] ),
    .I3(\soc.spi_video_ram_1.write_fifo.fifo_mem[15][20] ),
    .S0(_02713_),
    .S1(_02714_),
    .Z(_03578_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07937_ (.I(_02831_),
    .Z(_03579_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07938_ (.A1(_03577_),
    .A2(_03578_),
    .B(_03579_),
    .ZN(_03580_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _07939_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[0][20] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[1][20] ),
    .I2(\soc.spi_video_ram_1.write_fifo.fifo_mem[2][20] ),
    .I3(\soc.spi_video_ram_1.write_fifo.fifo_mem[3][20] ),
    .S0(_02764_),
    .S1(_02723_),
    .Z(_03581_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07940_ (.A1(_02768_),
    .A2(_03581_),
    .ZN(_03582_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _07941_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[4][20] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[5][20] ),
    .I2(\soc.spi_video_ram_1.write_fifo.fifo_mem[6][20] ),
    .I3(\soc.spi_video_ram_1.write_fifo.fifo_mem[7][20] ),
    .S0(_02764_),
    .S1(_02723_),
    .Z(_03583_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07942_ (.A1(_02571_),
    .A2(_03583_),
    .B(_02602_),
    .ZN(_03584_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _07943_ (.A1(_03576_),
    .A2(_03580_),
    .B1(_03582_),
    .B2(_03584_),
    .C(_02710_),
    .ZN(_03585_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _07944_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[24][20] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[25][20] ),
    .I2(\soc.spi_video_ram_1.write_fifo.fifo_mem[26][20] ),
    .I3(\soc.spi_video_ram_1.write_fifo.fifo_mem[27][20] ),
    .S0(_02713_),
    .S1(_02714_),
    .Z(_03586_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07945_ (.A1(_02678_),
    .A2(_03586_),
    .ZN(_03587_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _07946_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[28][20] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[29][20] ),
    .I2(\soc.spi_video_ram_1.write_fifo.fifo_mem[30][20] ),
    .I3(\soc.spi_video_ram_1.write_fifo.fifo_mem[31][20] ),
    .S0(_02713_),
    .S1(_02714_),
    .Z(_03588_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07947_ (.A1(_03577_),
    .A2(_03588_),
    .B(_03579_),
    .ZN(_03589_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _07948_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[16][20] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[17][20] ),
    .I2(\soc.spi_video_ram_1.write_fifo.fifo_mem[18][20] ),
    .I3(\soc.spi_video_ram_1.write_fifo.fifo_mem[19][20] ),
    .S0(_02764_),
    .S1(_02723_),
    .Z(_03590_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07949_ (.A1(_02768_),
    .A2(_03590_),
    .ZN(_03591_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _07950_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[20][20] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[21][20] ),
    .I2(\soc.spi_video_ram_1.write_fifo.fifo_mem[22][20] ),
    .I3(\soc.spi_video_ram_1.write_fifo.fifo_mem[23][20] ),
    .S0(_02769_),
    .S1(_02770_),
    .Z(_03592_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07951_ (.A1(_02571_),
    .A2(_03592_),
    .B(_02602_),
    .ZN(_03593_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _07952_ (.A1(_03587_),
    .A2(_03589_),
    .B1(_03591_),
    .B2(_03593_),
    .C(_02568_),
    .ZN(_03594_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07953_ (.A1(_03585_),
    .A2(_03594_),
    .ZN(_03595_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _07954_ (.A1(_02677_),
    .A2(_01392_),
    .A3(_02734_),
    .ZN(_03596_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07955_ (.A1(\soc.spi_video_ram_1.output_buffer[5] ),
    .A2(_02676_),
    .ZN(_03597_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07956_ (.A1(_03595_),
    .A2(_03596_),
    .B(_03597_),
    .ZN(_00251_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _07957_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[8][19] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[9][19] ),
    .I2(\soc.spi_video_ram_1.write_fifo.fifo_mem[10][19] ),
    .I3(\soc.spi_video_ram_1.write_fifo.fifo_mem[11][19] ),
    .S0(_02713_),
    .S1(_02737_),
    .Z(_03598_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07958_ (.A1(_02736_),
    .A2(_03598_),
    .ZN(_03599_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _07959_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[12][19] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[13][19] ),
    .I2(\soc.spi_video_ram_1.write_fifo.fifo_mem[14][19] ),
    .I3(\soc.spi_video_ram_1.write_fifo.fifo_mem[15][19] ),
    .S0(_02701_),
    .S1(_02737_),
    .Z(_03600_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07960_ (.A1(_03577_),
    .A2(_03600_),
    .B(_03579_),
    .ZN(_03601_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _07961_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[0][19] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[1][19] ),
    .I2(\soc.spi_video_ram_1.write_fifo.fifo_mem[2][19] ),
    .I3(\soc.spi_video_ram_1.write_fifo.fifo_mem[3][19] ),
    .S0(_02769_),
    .S1(_02770_),
    .Z(_03602_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07962_ (.A1(_02768_),
    .A2(_03602_),
    .ZN(_03603_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _07963_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[4][19] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[5][19] ),
    .I2(\soc.spi_video_ram_1.write_fifo.fifo_mem[6][19] ),
    .I3(\soc.spi_video_ram_1.write_fifo.fifo_mem[7][19] ),
    .S0(_02681_),
    .S1(_02758_),
    .Z(_03604_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07964_ (.A1(_02571_),
    .A2(_03604_),
    .B(_02602_),
    .ZN(_03605_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _07965_ (.A1(_03599_),
    .A2(_03601_),
    .B1(_03603_),
    .B2(_03605_),
    .C(_02710_),
    .ZN(_03606_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _07966_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[24][19] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[25][19] ),
    .I2(\soc.spi_video_ram_1.write_fifo.fifo_mem[26][19] ),
    .I3(\soc.spi_video_ram_1.write_fifo.fifo_mem[27][19] ),
    .S0(_02713_),
    .S1(_02737_),
    .Z(_03607_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07967_ (.A1(_02736_),
    .A2(_03607_),
    .ZN(_03608_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _07968_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[28][19] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[29][19] ),
    .I2(\soc.spi_video_ram_1.write_fifo.fifo_mem[30][19] ),
    .I3(\soc.spi_video_ram_1.write_fifo.fifo_mem[31][19] ),
    .S0(_02701_),
    .S1(_02737_),
    .Z(_03609_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07969_ (.A1(_03577_),
    .A2(_03609_),
    .B(_03579_),
    .ZN(_03610_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _07970_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[16][19] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[17][19] ),
    .I2(\soc.spi_video_ram_1.write_fifo.fifo_mem[18][19] ),
    .I3(\soc.spi_video_ram_1.write_fifo.fifo_mem[19][19] ),
    .S0(_02769_),
    .S1(_02770_),
    .Z(_03611_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07971_ (.A1(_02768_),
    .A2(_03611_),
    .ZN(_03612_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _07972_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[20][19] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[21][19] ),
    .I2(\soc.spi_video_ram_1.write_fifo.fifo_mem[22][19] ),
    .I3(\soc.spi_video_ram_1.write_fifo.fifo_mem[23][19] ),
    .S0(_02681_),
    .S1(_02758_),
    .Z(_03613_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07973_ (.A1(_02571_),
    .A2(_03613_),
    .B(_02602_),
    .ZN(_03614_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _07974_ (.A1(_03608_),
    .A2(_03610_),
    .B1(_03612_),
    .B2(_03614_),
    .C(_02568_),
    .ZN(_03615_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07975_ (.A1(_03606_),
    .A2(_03615_),
    .ZN(_03616_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _07976_ (.A1(_01539_),
    .A2(_02882_),
    .B1(_03596_),
    .B2(_03616_),
    .ZN(_00252_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _07977_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[8][18] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[9][18] ),
    .I2(\soc.spi_video_ram_1.write_fifo.fifo_mem[10][18] ),
    .I3(\soc.spi_video_ram_1.write_fifo.fifo_mem[11][18] ),
    .S0(_02701_),
    .S1(_02737_),
    .Z(_03617_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07978_ (.A1(_02736_),
    .A2(_03617_),
    .ZN(_03618_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _07979_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[12][18] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[13][18] ),
    .I2(\soc.spi_video_ram_1.write_fifo.fifo_mem[14][18] ),
    .I3(\soc.spi_video_ram_1.write_fifo.fifo_mem[15][18] ),
    .S0(_02726_),
    .S1(_03041_),
    .Z(_03619_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07980_ (.A1(_03577_),
    .A2(_03619_),
    .B(_03579_),
    .ZN(_03620_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _07981_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[0][18] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[1][18] ),
    .I2(\soc.spi_video_ram_1.write_fifo.fifo_mem[2][18] ),
    .I3(\soc.spi_video_ram_1.write_fifo.fifo_mem[3][18] ),
    .S0(_02681_),
    .S1(_02758_),
    .Z(_03621_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07982_ (.A1(_02768_),
    .A2(_03621_),
    .ZN(_03622_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _07983_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[4][18] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[5][18] ),
    .I2(\soc.spi_video_ram_1.write_fifo.fifo_mem[6][18] ),
    .I3(\soc.spi_video_ram_1.write_fifo.fifo_mem[7][18] ),
    .S0(_02717_),
    .S1(_02682_),
    .Z(_03623_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07984_ (.A1(_02685_),
    .A2(_03623_),
    .B(_02720_),
    .ZN(_03624_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _07985_ (.A1(_03618_),
    .A2(_03620_),
    .B1(_03622_),
    .B2(_03624_),
    .C(_02710_),
    .ZN(_03625_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _07986_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[16][18] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[17][18] ),
    .I2(\soc.spi_video_ram_1.write_fifo.fifo_mem[18][18] ),
    .I3(\soc.spi_video_ram_1.write_fifo.fifo_mem[19][18] ),
    .S0(_02701_),
    .S1(_03041_),
    .Z(_03626_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07987_ (.A1(_02736_),
    .A2(_03626_),
    .ZN(_03627_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _07988_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[20][18] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[21][18] ),
    .I2(\soc.spi_video_ram_1.write_fifo.fifo_mem[22][18] ),
    .I3(\soc.spi_video_ram_1.write_fifo.fifo_mem[23][18] ),
    .S0(_02726_),
    .S1(_03041_),
    .Z(_03628_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07989_ (.A1(_03577_),
    .A2(_03628_),
    .B(_02720_),
    .ZN(_03629_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _07990_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[24][18] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[25][18] ),
    .I2(\soc.spi_video_ram_1.write_fifo.fifo_mem[26][18] ),
    .I3(\soc.spi_video_ram_1.write_fifo.fifo_mem[27][18] ),
    .S0(_02681_),
    .S1(_02758_),
    .Z(_03630_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07991_ (.A1(_02678_),
    .A2(_03630_),
    .ZN(_03631_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _07992_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[28][18] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[29][18] ),
    .I2(\soc.spi_video_ram_1.write_fifo.fifo_mem[30][18] ),
    .I3(\soc.spi_video_ram_1.write_fifo.fifo_mem[31][18] ),
    .S0(_02717_),
    .S1(_02714_),
    .Z(_03632_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07993_ (.A1(_02685_),
    .A2(_03632_),
    .B(_03579_),
    .ZN(_03633_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _07994_ (.A1(_03627_),
    .A2(_03629_),
    .B1(_03631_),
    .B2(_03633_),
    .C(_02568_),
    .ZN(_03634_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07995_ (.A1(_03625_),
    .A2(_03634_),
    .ZN(_03635_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07996_ (.A1(\soc.spi_video_ram_1.output_buffer[3] ),
    .A2(_02676_),
    .ZN(_03636_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07997_ (.A1(_03596_),
    .A2(_03635_),
    .B(_03636_),
    .ZN(_00253_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _07998_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[8][17] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[9][17] ),
    .I2(\soc.spi_video_ram_1.write_fifo.fifo_mem[10][17] ),
    .I3(\soc.spi_video_ram_1.write_fifo.fifo_mem[11][17] ),
    .S0(_02701_),
    .S1(_02737_),
    .Z(_03637_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07999_ (.A1(_02736_),
    .A2(_03637_),
    .ZN(_03638_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _08000_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[12][17] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[13][17] ),
    .I2(\soc.spi_video_ram_1.write_fifo.fifo_mem[14][17] ),
    .I3(\soc.spi_video_ram_1.write_fifo.fifo_mem[15][17] ),
    .S0(_02726_),
    .S1(_03041_),
    .Z(_03639_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08001_ (.A1(_03577_),
    .A2(_03639_),
    .B(_03579_),
    .ZN(_03640_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _08002_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[0][17] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[1][17] ),
    .I2(\soc.spi_video_ram_1.write_fifo.fifo_mem[2][17] ),
    .I3(\soc.spi_video_ram_1.write_fifo.fifo_mem[3][17] ),
    .S0(_02769_),
    .S1(_02758_),
    .Z(_03641_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08003_ (.A1(_02768_),
    .A2(_03641_),
    .ZN(_03642_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _08004_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[4][17] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[5][17] ),
    .I2(\soc.spi_video_ram_1.write_fifo.fifo_mem[6][17] ),
    .I3(\soc.spi_video_ram_1.write_fifo.fifo_mem[7][17] ),
    .S0(_02717_),
    .S1(_02682_),
    .Z(_03643_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08005_ (.A1(_02685_),
    .A2(_03643_),
    .B(_02720_),
    .ZN(_03644_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _08006_ (.A1(_03638_),
    .A2(_03640_),
    .B1(_03642_),
    .B2(_03644_),
    .C(_02710_),
    .ZN(_03645_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _08007_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[24][17] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[25][17] ),
    .I2(\soc.spi_video_ram_1.write_fifo.fifo_mem[26][17] ),
    .I3(\soc.spi_video_ram_1.write_fifo.fifo_mem[27][17] ),
    .S0(_02701_),
    .S1(_02737_),
    .Z(_03646_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08008_ (.A1(_02736_),
    .A2(_03646_),
    .ZN(_03647_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _08009_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[28][17] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[29][17] ),
    .I2(\soc.spi_video_ram_1.write_fifo.fifo_mem[30][17] ),
    .I3(\soc.spi_video_ram_1.write_fifo.fifo_mem[31][17] ),
    .S0(_02726_),
    .S1(_03041_),
    .Z(_03648_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08010_ (.A1(_03577_),
    .A2(_03648_),
    .B(_03579_),
    .ZN(_03649_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _08011_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[16][17] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[17][17] ),
    .I2(\soc.spi_video_ram_1.write_fifo.fifo_mem[18][17] ),
    .I3(\soc.spi_video_ram_1.write_fifo.fifo_mem[19][17] ),
    .S0(_02681_),
    .S1(_02758_),
    .Z(_03650_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08012_ (.A1(_02678_),
    .A2(_03650_),
    .ZN(_03651_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _08013_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[20][17] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[21][17] ),
    .I2(\soc.spi_video_ram_1.write_fifo.fifo_mem[22][17] ),
    .I3(\soc.spi_video_ram_1.write_fifo.fifo_mem[23][17] ),
    .S0(_02717_),
    .S1(_02682_),
    .Z(_03652_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08014_ (.A1(_02685_),
    .A2(_03652_),
    .B(_02720_),
    .ZN(_03653_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _08015_ (.A1(_03647_),
    .A2(_03649_),
    .B1(_03651_),
    .B2(_03653_),
    .C(_02568_),
    .ZN(_03654_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08016_ (.A1(_03645_),
    .A2(_03654_),
    .ZN(_03655_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08017_ (.A1(\soc.spi_video_ram_1.output_buffer[2] ),
    .A2(_02675_),
    .ZN(_03656_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08018_ (.A1(_03596_),
    .A2(_03655_),
    .B(_03656_),
    .ZN(_00254_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _08019_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[0][16] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[1][16] ),
    .I2(\soc.spi_video_ram_1.write_fifo.fifo_mem[2][16] ),
    .I3(\soc.spi_video_ram_1.write_fifo.fifo_mem[3][16] ),
    .S0(_02701_),
    .S1(_02737_),
    .Z(_03657_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08020_ (.A1(_02736_),
    .A2(_03657_),
    .ZN(_03658_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _08021_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[4][16] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[5][16] ),
    .I2(\soc.spi_video_ram_1.write_fifo.fifo_mem[6][16] ),
    .I3(\soc.spi_video_ram_1.write_fifo.fifo_mem[7][16] ),
    .S0(_02701_),
    .S1(_03041_),
    .Z(_03659_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08022_ (.A1(_03577_),
    .A2(_03659_),
    .B(_02720_),
    .ZN(_03660_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _08023_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[8][16] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[9][16] ),
    .I2(\soc.spi_video_ram_1.write_fifo.fifo_mem[10][16] ),
    .I3(\soc.spi_video_ram_1.write_fifo.fifo_mem[11][16] ),
    .S0(_02769_),
    .S1(_02770_),
    .Z(_03661_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08024_ (.A1(_02768_),
    .A2(_03661_),
    .ZN(_03662_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _08025_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[12][16] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[13][16] ),
    .I2(\soc.spi_video_ram_1.write_fifo.fifo_mem[14][16] ),
    .I3(\soc.spi_video_ram_1.write_fifo.fifo_mem[15][16] ),
    .S0(_02717_),
    .S1(_02682_),
    .Z(_03663_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08026_ (.A1(_02685_),
    .A2(_03663_),
    .B(_03579_),
    .ZN(_03664_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _08027_ (.A1(_03658_),
    .A2(_03660_),
    .B1(_03662_),
    .B2(_03664_),
    .C(_02710_),
    .ZN(_03665_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _08028_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[24][16] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[25][16] ),
    .I2(\soc.spi_video_ram_1.write_fifo.fifo_mem[26][16] ),
    .I3(\soc.spi_video_ram_1.write_fifo.fifo_mem[27][16] ),
    .S0(_02701_),
    .S1(_02737_),
    .Z(_03666_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08029_ (.A1(_02736_),
    .A2(_03666_),
    .ZN(_03667_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _08030_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[28][16] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[29][16] ),
    .I2(\soc.spi_video_ram_1.write_fifo.fifo_mem[30][16] ),
    .I3(\soc.spi_video_ram_1.write_fifo.fifo_mem[31][16] ),
    .S0(_02726_),
    .S1(_03041_),
    .Z(_03668_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08031_ (.A1(_03577_),
    .A2(_03668_),
    .B(_03579_),
    .ZN(_03669_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _08032_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[16][16] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[17][16] ),
    .I2(\soc.spi_video_ram_1.write_fifo.fifo_mem[18][16] ),
    .I3(\soc.spi_video_ram_1.write_fifo.fifo_mem[19][16] ),
    .S0(_02681_),
    .S1(_02758_),
    .Z(_03670_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08033_ (.A1(_02768_),
    .A2(_03670_),
    .ZN(_03671_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _08034_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[20][16] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[21][16] ),
    .I2(\soc.spi_video_ram_1.write_fifo.fifo_mem[22][16] ),
    .I3(\soc.spi_video_ram_1.write_fifo.fifo_mem[23][16] ),
    .S0(_02717_),
    .S1(_02682_),
    .Z(_03672_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08035_ (.A1(_02685_),
    .A2(_03672_),
    .B(_02720_),
    .ZN(_03673_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _08036_ (.A1(_03667_),
    .A2(_03669_),
    .B1(_03671_),
    .B2(_03673_),
    .C(_02568_),
    .ZN(_03674_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08037_ (.A1(_03665_),
    .A2(_03674_),
    .ZN(_03675_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08038_ (.A1(\soc.spi_video_ram_1.output_buffer[1] ),
    .A2(_02675_),
    .ZN(_03676_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08039_ (.A1(_03596_),
    .A2(_03675_),
    .B(_03676_),
    .ZN(_00255_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08040_ (.A1(_02115_),
    .A2(_01403_),
    .ZN(_03677_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _08041_ (.A1(_02116_),
    .A2(_01441_),
    .A3(_03677_),
    .ZN(_03678_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _08042_ (.I(_03678_),
    .Z(_03679_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _08043_ (.I(_03679_),
    .Z(_03680_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08044_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[11][0] ),
    .I1(_02310_),
    .S(_03680_),
    .Z(_03681_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08045_ (.I(_03681_),
    .Z(_00256_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08046_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[11][1] ),
    .I1(_02393_),
    .S(_03680_),
    .Z(_03682_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08047_ (.I(_03682_),
    .Z(_00257_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08048_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[11][2] ),
    .I1(_02395_),
    .S(_03680_),
    .Z(_03683_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08049_ (.I(_03683_),
    .Z(_00258_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08050_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[11][3] ),
    .I1(_02397_),
    .S(_03680_),
    .Z(_03684_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08051_ (.I(_03684_),
    .Z(_00259_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08052_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[11][4] ),
    .I1(_02399_),
    .S(_03680_),
    .Z(_03685_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08053_ (.I(_03685_),
    .Z(_00260_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08054_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[11][5] ),
    .I1(_02401_),
    .S(_03680_),
    .Z(_03686_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08055_ (.I(_03686_),
    .Z(_00261_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08056_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[11][6] ),
    .I1(_02403_),
    .S(_03680_),
    .Z(_03687_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08057_ (.I(_03687_),
    .Z(_00262_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08058_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[11][7] ),
    .I1(_02405_),
    .S(_03680_),
    .Z(_03688_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08059_ (.I(_03688_),
    .Z(_00263_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08060_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[11][8] ),
    .I1(_02407_),
    .S(_03680_),
    .Z(_03689_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08061_ (.I(_03689_),
    .Z(_00264_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08062_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[11][9] ),
    .I1(_02409_),
    .S(_03680_),
    .Z(_03690_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08063_ (.I(_03690_),
    .Z(_00265_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _08064_ (.I(_03678_),
    .Z(_03691_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08065_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[11][10] ),
    .I1(_02411_),
    .S(_03691_),
    .Z(_03692_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08066_ (.I(_03692_),
    .Z(_00266_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08067_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[11][11] ),
    .I1(_02414_),
    .S(_03691_),
    .Z(_03693_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08068_ (.I(_03693_),
    .Z(_00267_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08069_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[11][12] ),
    .I1(_02242_),
    .S(_03691_),
    .Z(_03694_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08070_ (.I(_03694_),
    .Z(_00268_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08071_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[11][13] ),
    .I1(_02244_),
    .S(_03691_),
    .Z(_03695_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08072_ (.I(_03695_),
    .Z(_00269_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08073_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[11][14] ),
    .I1(_02246_),
    .S(_03691_),
    .Z(_03696_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08074_ (.I(_03696_),
    .Z(_00270_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08075_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[11][15] ),
    .I1(_02248_),
    .S(_03691_),
    .Z(_03697_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08076_ (.I(_03697_),
    .Z(_00271_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08077_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[11][16] ),
    .I1(_02335_),
    .S(_03691_),
    .Z(_03698_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08078_ (.I(_03698_),
    .Z(_00272_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08079_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[11][17] ),
    .I1(_02337_),
    .S(_03691_),
    .Z(_03699_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08080_ (.I(_03699_),
    .Z(_00273_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08081_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[11][18] ),
    .I1(_02339_),
    .S(_03691_),
    .Z(_03700_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08082_ (.I(_03700_),
    .Z(_00274_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08083_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[11][19] ),
    .I1(_02341_),
    .S(_03691_),
    .Z(_03701_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08084_ (.I(_03701_),
    .Z(_00275_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08085_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[11][20] ),
    .I1(_02343_),
    .S(_03679_),
    .Z(_03702_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08086_ (.I(_03702_),
    .Z(_00276_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08087_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[11][21] ),
    .I1(_02260_),
    .S(_03679_),
    .Z(_03703_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08088_ (.I(_03703_),
    .Z(_00277_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08089_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[11][22] ),
    .I1(_02262_),
    .S(_03679_),
    .Z(_03704_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08090_ (.I(_03704_),
    .Z(_00278_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08091_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[11][23] ),
    .I1(_02264_),
    .S(_03679_),
    .Z(_03705_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08092_ (.I(_03705_),
    .Z(_00279_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08093_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[11][24] ),
    .I1(_02266_),
    .S(_03679_),
    .Z(_03706_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08094_ (.I(_03706_),
    .Z(_00280_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08095_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[11][25] ),
    .I1(_02268_),
    .S(_03679_),
    .Z(_03707_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08096_ (.I(_03707_),
    .Z(_00281_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08097_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[11][26] ),
    .I1(_02270_),
    .S(_03679_),
    .Z(_03708_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08098_ (.I(_03708_),
    .Z(_00282_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08099_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[11][27] ),
    .I1(_02351_),
    .S(_03679_),
    .Z(_03709_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08100_ (.I(_03709_),
    .Z(_00283_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08101_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[11][28] ),
    .I1(_02353_),
    .S(_03679_),
    .Z(_03710_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08102_ (.I(_03710_),
    .Z(_00284_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _08103_ (.A1(\soc.video_generator_1.h_count[4] ),
    .A2(\soc.video_generator_1.h_count[7] ),
    .A3(\soc.video_generator_1.h_count[6] ),
    .ZN(_03711_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _08104_ (.A1(_01836_),
    .A2(_01968_),
    .A3(_01993_),
    .A4(_03711_),
    .ZN(_03712_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _08105_ (.A1(_01959_),
    .A2(_03712_),
    .B(_01380_),
    .ZN(_03713_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08106_ (.A1(\soc.display_clks_before_active[0] ),
    .A2(_03713_),
    .ZN(_00285_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08107_ (.I(_01395_),
    .Z(_03714_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08108_ (.A1(_01926_),
    .A2(_01994_),
    .ZN(_03715_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _08109_ (.A1(_03714_),
    .A2(_01968_),
    .A3(_03715_),
    .ZN(_00286_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08110_ (.A1(\soc.video_generator_1.h_count[2] ),
    .A2(_01990_),
    .Z(_03716_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08111_ (.A1(_03713_),
    .A2(_03716_),
    .ZN(_00287_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _08112_ (.A1(\soc.video_generator_1.h_count[3] ),
    .A2(\soc.video_generator_1.h_count[2] ),
    .A3(_03715_),
    .Z(_03717_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08113_ (.A1(\soc.video_generator_1.h_count[2] ),
    .A2(_03715_),
    .B(\soc.video_generator_1.h_count[3] ),
    .ZN(_03718_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _08114_ (.A1(_03713_),
    .A2(_03717_),
    .A3(_03718_),
    .ZN(_00288_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _08115_ (.A1(\soc.video_generator_1.h_count[4] ),
    .A2(_03717_),
    .Z(_03719_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08116_ (.A1(\soc.video_generator_1.h_count[4] ),
    .A2(_03717_),
    .ZN(_03720_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _08117_ (.A1(_03713_),
    .A2(_03719_),
    .A3(_03720_),
    .ZN(_00289_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _08118_ (.A1(_01836_),
    .A2(_03719_),
    .ZN(_03721_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08119_ (.A1(_03713_),
    .A2(_03721_),
    .ZN(_00290_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08120_ (.A1(_01836_),
    .A2(_03719_),
    .B(\soc.video_generator_1.h_count[6] ),
    .ZN(_03722_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _08121_ (.A1(_01836_),
    .A2(\soc.video_generator_1.h_count[6] ),
    .A3(_03719_),
    .Z(_03723_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _08122_ (.A1(_03713_),
    .A2(_03722_),
    .A3(_03723_),
    .ZN(_00291_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08123_ (.A1(\soc.video_generator_1.h_count[7] ),
    .A2(_03723_),
    .ZN(_03724_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _08124_ (.A1(\soc.video_generator_1.h_count[7] ),
    .A2(_03723_),
    .Z(_03725_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _08125_ (.A1(_03713_),
    .A2(_03724_),
    .A3(_03725_),
    .ZN(_00292_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _08126_ (.A1(_01959_),
    .A2(_03712_),
    .B1(_03725_),
    .B2(\soc.video_generator_1.h_count[8] ),
    .C(_01380_),
    .ZN(_03726_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08127_ (.A1(\soc.video_generator_1.h_count[8] ),
    .A2(_03725_),
    .B(_03726_),
    .ZN(_00293_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08128_ (.A1(\soc.video_generator_1.h_count[8] ),
    .A2(_03725_),
    .ZN(_03727_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _08129_ (.A1(\soc.video_generator_1.h_count[9] ),
    .A2(_03727_),
    .Z(_03728_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08130_ (.A1(_03713_),
    .A2(_03728_),
    .ZN(_00294_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08131_ (.A1(_02116_),
    .A2(_03677_),
    .ZN(_03729_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08132_ (.A1(_02114_),
    .A2(_03729_),
    .ZN(_03730_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _08133_ (.I(_03730_),
    .Z(_03731_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _08134_ (.I(_03731_),
    .Z(_03732_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08135_ (.I0(_02113_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[10][0] ),
    .S(_03732_),
    .Z(_03733_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08136_ (.I(_03733_),
    .Z(_00295_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08137_ (.I0(_02122_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[10][1] ),
    .S(_03732_),
    .Z(_03734_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08138_ (.I(_03734_),
    .Z(_00296_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08139_ (.I0(_02124_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[10][2] ),
    .S(_03732_),
    .Z(_03735_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08140_ (.I(_03735_),
    .Z(_00297_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08141_ (.I0(_02126_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[10][3] ),
    .S(_03732_),
    .Z(_03736_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08142_ (.I(_03736_),
    .Z(_00298_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08143_ (.I0(_02128_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[10][4] ),
    .S(_03732_),
    .Z(_03737_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08144_ (.I(_03737_),
    .Z(_00299_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08145_ (.I0(_02130_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[10][5] ),
    .S(_03732_),
    .Z(_03738_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08146_ (.I(_03738_),
    .Z(_00300_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08147_ (.I0(_02132_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[10][6] ),
    .S(_03732_),
    .Z(_03739_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08148_ (.I(_03739_),
    .Z(_00301_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08149_ (.I0(_02134_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[10][7] ),
    .S(_03732_),
    .Z(_03740_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08150_ (.I(_03740_),
    .Z(_00302_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08151_ (.I0(_02136_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[10][8] ),
    .S(_03732_),
    .Z(_03741_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08152_ (.I(_03741_),
    .Z(_00303_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08153_ (.I0(_02138_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[10][9] ),
    .S(_03732_),
    .Z(_03742_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08154_ (.I(_03742_),
    .Z(_00304_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _08155_ (.I(_03730_),
    .Z(_03743_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08156_ (.I0(_02140_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[10][10] ),
    .S(_03743_),
    .Z(_03744_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08157_ (.I(_03744_),
    .Z(_00305_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08158_ (.I0(_02143_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[10][11] ),
    .S(_03743_),
    .Z(_03745_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08159_ (.I(_03745_),
    .Z(_00306_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08160_ (.I0(_02145_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[10][12] ),
    .S(_03743_),
    .Z(_03746_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08161_ (.I(_03746_),
    .Z(_00307_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08162_ (.I0(_02147_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[10][13] ),
    .S(_03743_),
    .Z(_03747_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08163_ (.I(_03747_),
    .Z(_00308_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08164_ (.I0(_02149_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[10][14] ),
    .S(_03743_),
    .Z(_03748_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08165_ (.I(_03748_),
    .Z(_00309_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08166_ (.I0(_02151_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[10][15] ),
    .S(_03743_),
    .Z(_03749_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08167_ (.I(_03749_),
    .Z(_00310_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08168_ (.I0(_02153_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[10][16] ),
    .S(_03743_),
    .Z(_03750_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08169_ (.I(_03750_),
    .Z(_00311_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08170_ (.I0(_02155_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[10][17] ),
    .S(_03743_),
    .Z(_03751_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08171_ (.I(_03751_),
    .Z(_00312_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08172_ (.I0(_02157_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[10][18] ),
    .S(_03743_),
    .Z(_03752_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08173_ (.I(_03752_),
    .Z(_00313_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08174_ (.I0(_02159_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[10][19] ),
    .S(_03743_),
    .Z(_03753_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08175_ (.I(_03753_),
    .Z(_00314_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08176_ (.I0(_02161_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[10][20] ),
    .S(_03731_),
    .Z(_03754_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08177_ (.I(_03754_),
    .Z(_00315_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08178_ (.I0(_02163_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[10][21] ),
    .S(_03731_),
    .Z(_03755_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08179_ (.I(_03755_),
    .Z(_00316_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08180_ (.I0(_02165_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[10][22] ),
    .S(_03731_),
    .Z(_03756_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08181_ (.I(_03756_),
    .Z(_00317_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08182_ (.I0(_02167_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[10][23] ),
    .S(_03731_),
    .Z(_03757_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08183_ (.I(_03757_),
    .Z(_00318_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08184_ (.I0(_02169_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[10][24] ),
    .S(_03731_),
    .Z(_03758_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08185_ (.I(_03758_),
    .Z(_00319_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08186_ (.I0(_02171_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[10][25] ),
    .S(_03731_),
    .Z(_03759_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08187_ (.I(_03759_),
    .Z(_00320_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08188_ (.I0(_02173_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[10][26] ),
    .S(_03731_),
    .Z(_03760_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08189_ (.I(_03760_),
    .Z(_00321_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08190_ (.I0(_02175_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[10][27] ),
    .S(_03731_),
    .Z(_03761_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08191_ (.I(_03761_),
    .Z(_00322_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08192_ (.I0(_02177_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[10][28] ),
    .S(_03731_),
    .Z(_03762_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08193_ (.I(_03762_),
    .Z(_00323_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08194_ (.A1(_02433_),
    .A2(_02437_),
    .ZN(_03763_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08195_ (.A1(_03763_),
    .A2(_02458_),
    .ZN(_03764_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _08196_ (.A1(_02442_),
    .A2(_02463_),
    .ZN(_03765_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08197_ (.A1(_02445_),
    .A2(_03765_),
    .ZN(_03766_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _08198_ (.A1(_02443_),
    .A2(_02463_),
    .ZN(_03767_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08199_ (.A1(\soc.rom_encoder_0.output_buffer[16] ),
    .A2(_03766_),
    .B1(_03767_),
    .B2(\soc.rom_encoder_0.request_data_out[12] ),
    .ZN(_03768_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08200_ (.A1(_02460_),
    .A2(_03764_),
    .ZN(_03769_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08201_ (.I(\soc.rom_encoder_0.output_buffer[16] ),
    .ZN(_03770_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08202_ (.A1(_03764_),
    .A2(_03768_),
    .B1(_03769_),
    .B2(_03770_),
    .ZN(_03771_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08203_ (.A1(\soc.rom_encoder_0.initializing_step[1] ),
    .A2(_02459_),
    .B(\soc.rom_encoder_0.initializing_step[2] ),
    .ZN(_03772_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _08204_ (.A1(\soc.rom_encoder_0.initializing_step[4] ),
    .A2(\soc.rom_encoder_0.initializing_step[3] ),
    .A3(_03772_),
    .ZN(_03773_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _08205_ (.A1(_03763_),
    .A2(_02449_),
    .A3(_03773_),
    .ZN(_03774_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _08206_ (.A1(\soc.rom_encoder_0.initializing_step[4] ),
    .A2(\soc.rom_encoder_0.initializing_step[3] ),
    .A3(_02452_),
    .ZN(_03775_));
 gf180mcu_fd_sc_mcu7t5v0__oai33_1 _08207_ (.A1(_02452_),
    .A2(_03771_),
    .A3(_03774_),
    .B1(_03775_),
    .B2(_02540_),
    .B3(net64),
    .ZN(_03776_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08208_ (.A1(_01381_),
    .A2(_03776_),
    .ZN(_00324_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08209_ (.A1(\soc.ram_encoder_0.initializing_step[0] ),
    .A2(_02550_),
    .ZN(_03777_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _08210_ (.A1(_02484_),
    .A2(_02491_),
    .A3(_02479_),
    .ZN(_03778_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08211_ (.I(_03778_),
    .ZN(_03779_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08212_ (.A1(_02493_),
    .A2(_03777_),
    .B(_03779_),
    .C(_02487_),
    .ZN(_03780_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08213_ (.I(_03780_),
    .Z(_03781_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08214_ (.A1(\soc.ram_encoder_0.request_address[4] ),
    .A2(_02506_),
    .B1(_03781_),
    .B2(\soc.ram_encoder_0.output_buffer[1] ),
    .ZN(_03782_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08215_ (.A1(\soc.ram_encoder_0.output_buffer[5] ),
    .A2(_02563_),
    .ZN(_03783_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08216_ (.A1(_02556_),
    .A2(_03782_),
    .B(_03783_),
    .ZN(_00325_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08217_ (.A1(\soc.ram_encoder_0.request_address[5] ),
    .A2(_02506_),
    .B1(_03781_),
    .B2(\soc.ram_encoder_0.output_buffer[2] ),
    .ZN(_03784_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08218_ (.A1(\soc.ram_encoder_0.output_buffer[6] ),
    .A2(_02563_),
    .ZN(_03785_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08219_ (.A1(_02556_),
    .A2(_03784_),
    .B(_03785_),
    .ZN(_00326_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08220_ (.A1(\soc.ram_encoder_0.request_address[6] ),
    .A2(_02506_),
    .B1(_03781_),
    .B2(\soc.ram_encoder_0.output_buffer[3] ),
    .ZN(_03786_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08221_ (.A1(\soc.ram_encoder_0.output_buffer[7] ),
    .A2(_02563_),
    .ZN(_03787_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08222_ (.A1(_02556_),
    .A2(_03786_),
    .B(_03787_),
    .ZN(_00327_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _08223_ (.A1(_02503_),
    .A2(_02483_),
    .ZN(_03788_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08224_ (.I(_03788_),
    .Z(_03789_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _08225_ (.A1(\soc.ram_encoder_0.request_address[7] ),
    .A2(_02506_),
    .Z(_03790_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _08226_ (.A1(\soc.ram_encoder_0.output_buffer[4] ),
    .A2(_03781_),
    .B1(_03789_),
    .B2(\soc.ram_encoder_0.request_data_out[0] ),
    .C(_03790_),
    .ZN(_03791_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08227_ (.A1(\soc.ram_encoder_0.output_buffer[8] ),
    .A2(_02563_),
    .ZN(_03792_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08228_ (.A1(_02556_),
    .A2(_03791_),
    .B(_03792_),
    .ZN(_00328_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _08229_ (.A1(\soc.ram_encoder_0.request_address[8] ),
    .A2(_02505_),
    .Z(_03793_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _08230_ (.A1(\soc.ram_encoder_0.output_buffer[5] ),
    .A2(_03781_),
    .B1(_03789_),
    .B2(\soc.ram_encoder_0.request_data_out[1] ),
    .C(_03793_),
    .ZN(_03794_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08231_ (.A1(\soc.ram_encoder_0.output_buffer[9] ),
    .A2(_02563_),
    .ZN(_03795_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08232_ (.A1(_02556_),
    .A2(_03794_),
    .B(_03795_),
    .ZN(_00329_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _08233_ (.A1(\soc.ram_encoder_0.request_address[9] ),
    .A2(_02505_),
    .Z(_03796_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _08234_ (.A1(\soc.ram_encoder_0.output_buffer[6] ),
    .A2(_03781_),
    .B1(_03789_),
    .B2(\soc.ram_encoder_0.request_data_out[2] ),
    .C(_03796_),
    .ZN(_03797_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08235_ (.A1(\soc.ram_encoder_0.output_buffer[10] ),
    .A2(_02563_),
    .ZN(_03798_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08236_ (.A1(_02556_),
    .A2(_03797_),
    .B(_03798_),
    .ZN(_00330_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _08237_ (.A1(\soc.ram_encoder_0.request_address[10] ),
    .A2(_02505_),
    .Z(_03799_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _08238_ (.A1(\soc.ram_encoder_0.output_buffer[7] ),
    .A2(_03781_),
    .B1(_03789_),
    .B2(\soc.ram_encoder_0.request_data_out[3] ),
    .C(_03799_),
    .ZN(_03800_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08239_ (.A1(\soc.ram_encoder_0.output_buffer[11] ),
    .A2(_02563_),
    .ZN(_03801_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08240_ (.A1(_02558_),
    .A2(_03800_),
    .B(_03801_),
    .ZN(_00331_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _08241_ (.A1(\soc.ram_encoder_0.request_address[11] ),
    .A2(_02505_),
    .Z(_03802_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _08242_ (.A1(\soc.ram_encoder_0.output_buffer[8] ),
    .A2(_03781_),
    .B1(_03789_),
    .B2(\soc.ram_encoder_0.request_data_out[4] ),
    .C(_03802_),
    .ZN(_03803_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08243_ (.A1(\soc.ram_encoder_0.output_buffer[12] ),
    .A2(_02563_),
    .ZN(_03804_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08244_ (.A1(_02558_),
    .A2(_03803_),
    .B(_03804_),
    .ZN(_00332_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _08245_ (.A1(\soc.ram_encoder_0.request_address[12] ),
    .A2(_02505_),
    .Z(_03805_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _08246_ (.A1(\soc.ram_encoder_0.output_buffer[9] ),
    .A2(_03781_),
    .B1(_03789_),
    .B2(\soc.ram_encoder_0.request_data_out[5] ),
    .C(_03805_),
    .ZN(_03806_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08247_ (.A1(\soc.ram_encoder_0.output_buffer[13] ),
    .A2(_02555_),
    .ZN(_03807_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08248_ (.A1(_02558_),
    .A2(_03806_),
    .B(_03807_),
    .ZN(_00333_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _08249_ (.A1(\soc.ram_encoder_0.request_address[13] ),
    .A2(_02505_),
    .Z(_03808_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _08250_ (.A1(\soc.ram_encoder_0.output_buffer[10] ),
    .A2(_03781_),
    .B1(_03789_),
    .B2(\soc.ram_encoder_0.request_data_out[6] ),
    .C(_03808_),
    .ZN(_03809_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08251_ (.A1(\soc.ram_encoder_0.output_buffer[14] ),
    .A2(_02555_),
    .ZN(_03810_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08252_ (.A1(_02558_),
    .A2(_03809_),
    .B(_03810_),
    .ZN(_00334_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _08253_ (.A1(\soc.ram_encoder_0.output_buffer[11] ),
    .A2(_03780_),
    .Z(_03811_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _08254_ (.A1(\soc.ram_encoder_0.request_address[14] ),
    .A2(_02506_),
    .B1(_03789_),
    .B2(\soc.ram_encoder_0.request_data_out[7] ),
    .C(_03811_),
    .ZN(_03812_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08255_ (.A1(\soc.ram_encoder_0.output_buffer[15] ),
    .A2(_02555_),
    .ZN(_03813_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08256_ (.A1(_02558_),
    .A2(_03812_),
    .B(_03813_),
    .ZN(_00335_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _08257_ (.A1(_02480_),
    .A2(_02498_),
    .A3(_03779_),
    .ZN(_03814_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08258_ (.A1(\soc.ram_encoder_0.output_buffer[12] ),
    .A2(_03814_),
    .ZN(_03815_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08259_ (.I(\soc.ram_encoder_0.request_write ),
    .ZN(_03816_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _08260_ (.A1(_02500_),
    .A2(_03777_),
    .Z(_03817_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _08261_ (.A1(_03816_),
    .A2(_02510_),
    .B1(_03788_),
    .B2(\soc.ram_encoder_0.request_data_out[8] ),
    .C(_03817_),
    .ZN(_03818_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08262_ (.A1(_03815_),
    .A2(_03818_),
    .ZN(_03819_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08263_ (.I0(_03819_),
    .I1(\soc.ram_encoder_0.output_buffer[16] ),
    .S(_02555_),
    .Z(_03820_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08264_ (.I(_03820_),
    .Z(_00336_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08265_ (.A1(_02479_),
    .A2(_02493_),
    .ZN(_03821_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _08266_ (.A1(\soc.ram_encoder_0.output_buffer[13] ),
    .A2(_03817_),
    .Z(_03822_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _08267_ (.A1(\soc.ram_encoder_0.request_data_out[9] ),
    .A2(_03789_),
    .B1(_03821_),
    .B2(_03822_),
    .C(_02510_),
    .ZN(_03823_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08268_ (.A1(\soc.ram_encoder_0.output_buffer[17] ),
    .A2(_02555_),
    .ZN(_03824_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08269_ (.A1(_02558_),
    .A2(_03823_),
    .B(_03824_),
    .ZN(_00337_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _08270_ (.A1(\soc.ram_encoder_0.output_buffer[14] ),
    .A2(_03814_),
    .B1(_03789_),
    .B2(\soc.ram_encoder_0.request_data_out[10] ),
    .C(_03817_),
    .ZN(_03825_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08271_ (.A1(\soc.ram_encoder_0.output_buffer[18] ),
    .A2(_02555_),
    .ZN(_03826_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08272_ (.A1(_02558_),
    .A2(_03825_),
    .B(_03826_),
    .ZN(_00338_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _08273_ (.A1(\soc.ram_encoder_0.output_buffer[15] ),
    .A2(_03814_),
    .B1(_03788_),
    .B2(\soc.ram_encoder_0.request_data_out[11] ),
    .C(_03817_),
    .ZN(_03827_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08274_ (.A1(\soc.ram_encoder_0.output_buffer[19] ),
    .A2(_02555_),
    .ZN(_03828_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08275_ (.A1(_02558_),
    .A2(_03827_),
    .B(_03828_),
    .ZN(_00339_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08276_ (.A1(_02179_),
    .A2(_02276_),
    .ZN(_03829_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _08277_ (.I(_03829_),
    .Z(_03830_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _08278_ (.I(_03830_),
    .Z(_03831_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08279_ (.I0(_02113_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[1][0] ),
    .S(_03831_),
    .Z(_03832_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08280_ (.I(_03832_),
    .Z(_00340_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08281_ (.I0(_02122_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[1][1] ),
    .S(_03831_),
    .Z(_03833_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08282_ (.I(_03833_),
    .Z(_00341_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08283_ (.I0(_02124_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[1][2] ),
    .S(_03831_),
    .Z(_03834_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08284_ (.I(_03834_),
    .Z(_00342_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08285_ (.I0(_02126_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[1][3] ),
    .S(_03831_),
    .Z(_03835_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08286_ (.I(_03835_),
    .Z(_00343_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08287_ (.I0(_02128_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[1][4] ),
    .S(_03831_),
    .Z(_03836_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08288_ (.I(_03836_),
    .Z(_00344_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08289_ (.I0(_02130_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[1][5] ),
    .S(_03831_),
    .Z(_03837_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08290_ (.I(_03837_),
    .Z(_00345_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08291_ (.I0(_02132_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[1][6] ),
    .S(_03831_),
    .Z(_03838_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08292_ (.I(_03838_),
    .Z(_00346_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08293_ (.I0(_02134_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[1][7] ),
    .S(_03831_),
    .Z(_03839_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08294_ (.I(_03839_),
    .Z(_00347_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08295_ (.I0(_02136_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[1][8] ),
    .S(_03831_),
    .Z(_03840_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08296_ (.I(_03840_),
    .Z(_00348_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08297_ (.I0(_02138_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[1][9] ),
    .S(_03831_),
    .Z(_03841_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08298_ (.I(_03841_),
    .Z(_00349_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _08299_ (.I(_03829_),
    .Z(_03842_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08300_ (.I0(_02140_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[1][10] ),
    .S(_03842_),
    .Z(_03843_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08301_ (.I(_03843_),
    .Z(_00350_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08302_ (.I0(_02143_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[1][11] ),
    .S(_03842_),
    .Z(_03844_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08303_ (.I(_03844_),
    .Z(_00351_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08304_ (.I0(_02145_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[1][12] ),
    .S(_03842_),
    .Z(_03845_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08305_ (.I(_03845_),
    .Z(_00352_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08306_ (.I0(_02147_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[1][13] ),
    .S(_03842_),
    .Z(_03846_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08307_ (.I(_03846_),
    .Z(_00353_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08308_ (.I0(_02149_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[1][14] ),
    .S(_03842_),
    .Z(_03847_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08309_ (.I(_03847_),
    .Z(_00354_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08310_ (.I0(_02151_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[1][15] ),
    .S(_03842_),
    .Z(_03848_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08311_ (.I(_03848_),
    .Z(_00355_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08312_ (.I0(_02153_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[1][16] ),
    .S(_03842_),
    .Z(_03849_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08313_ (.I(_03849_),
    .Z(_00356_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08314_ (.I0(_02155_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[1][17] ),
    .S(_03842_),
    .Z(_03850_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08315_ (.I(_03850_),
    .Z(_00357_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08316_ (.I0(_02157_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[1][18] ),
    .S(_03842_),
    .Z(_03851_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08317_ (.I(_03851_),
    .Z(_00358_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08318_ (.I0(_02159_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[1][19] ),
    .S(_03842_),
    .Z(_03852_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08319_ (.I(_03852_),
    .Z(_00359_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08320_ (.I0(_02161_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[1][20] ),
    .S(_03830_),
    .Z(_03853_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08321_ (.I(_03853_),
    .Z(_00360_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08322_ (.I0(_02163_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[1][21] ),
    .S(_03830_),
    .Z(_03854_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08323_ (.I(_03854_),
    .Z(_00361_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08324_ (.I0(_02165_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[1][22] ),
    .S(_03830_),
    .Z(_03855_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08325_ (.I(_03855_),
    .Z(_00362_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08326_ (.I0(_02167_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[1][23] ),
    .S(_03830_),
    .Z(_03856_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08327_ (.I(_03856_),
    .Z(_00363_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08328_ (.I0(_02169_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[1][24] ),
    .S(_03830_),
    .Z(_03857_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08329_ (.I(_03857_),
    .Z(_00364_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08330_ (.I0(_02171_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[1][25] ),
    .S(_03830_),
    .Z(_03858_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08331_ (.I(_03858_),
    .Z(_00365_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08332_ (.I0(_02173_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[1][26] ),
    .S(_03830_),
    .Z(_03859_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08333_ (.I(_03859_),
    .Z(_00366_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08334_ (.I0(_02175_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[1][27] ),
    .S(_03830_),
    .Z(_03860_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08335_ (.I(_03860_),
    .Z(_00367_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08336_ (.I0(_02177_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[1][28] ),
    .S(_03830_),
    .Z(_03861_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08337_ (.I(_03861_),
    .Z(_00368_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _08338_ (.I(\soc.spi_video_ram_1.write_fifo.write_pointer[2] ),
    .ZN(_03862_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _08339_ (.A1(\soc.spi_video_ram_1.write_fifo.write_pointer[4] ),
    .A2(_01403_),
    .A3(_03862_),
    .ZN(_03863_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08340_ (.A1(_02388_),
    .A2(_03863_),
    .ZN(_03864_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _08341_ (.I(_03864_),
    .Z(_03865_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _08342_ (.I(_03865_),
    .Z(_03866_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08343_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[26][0] ),
    .I1(_02310_),
    .S(_03866_),
    .Z(_03867_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08344_ (.I(_03867_),
    .Z(_00369_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08345_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[26][1] ),
    .I1(_02393_),
    .S(_03866_),
    .Z(_03868_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08346_ (.I(_03868_),
    .Z(_00370_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08347_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[26][2] ),
    .I1(_02395_),
    .S(_03866_),
    .Z(_03869_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08348_ (.I(_03869_),
    .Z(_00371_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08349_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[26][3] ),
    .I1(_02397_),
    .S(_03866_),
    .Z(_03870_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08350_ (.I(_03870_),
    .Z(_00372_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08351_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[26][4] ),
    .I1(_02399_),
    .S(_03866_),
    .Z(_03871_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08352_ (.I(_03871_),
    .Z(_00373_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08353_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[26][5] ),
    .I1(_02401_),
    .S(_03866_),
    .Z(_03872_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08354_ (.I(_03872_),
    .Z(_00374_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08355_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[26][6] ),
    .I1(_02403_),
    .S(_03866_),
    .Z(_03873_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08356_ (.I(_03873_),
    .Z(_00375_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08357_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[26][7] ),
    .I1(_02405_),
    .S(_03866_),
    .Z(_03874_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08358_ (.I(_03874_),
    .Z(_00376_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08359_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[26][8] ),
    .I1(_02407_),
    .S(_03866_),
    .Z(_03875_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08360_ (.I(_03875_),
    .Z(_00377_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08361_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[26][9] ),
    .I1(_02409_),
    .S(_03866_),
    .Z(_03876_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08362_ (.I(_03876_),
    .Z(_00378_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _08363_ (.I(_03864_),
    .Z(_03877_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08364_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[26][10] ),
    .I1(_02411_),
    .S(_03877_),
    .Z(_03878_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08365_ (.I(_03878_),
    .Z(_00379_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08366_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[26][11] ),
    .I1(_02414_),
    .S(_03877_),
    .Z(_03879_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08367_ (.I(_03879_),
    .Z(_00380_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08368_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[26][12] ),
    .I1(_02242_),
    .S(_03877_),
    .Z(_03880_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08369_ (.I(_03880_),
    .Z(_00381_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08370_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[26][13] ),
    .I1(_02244_),
    .S(_03877_),
    .Z(_03881_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08371_ (.I(_03881_),
    .Z(_00382_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08372_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[26][14] ),
    .I1(_02246_),
    .S(_03877_),
    .Z(_03882_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08373_ (.I(_03882_),
    .Z(_00383_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08374_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[26][15] ),
    .I1(_02248_),
    .S(_03877_),
    .Z(_03883_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08375_ (.I(_03883_),
    .Z(_00384_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08376_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[26][16] ),
    .I1(_02335_),
    .S(_03877_),
    .Z(_03884_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08377_ (.I(_03884_),
    .Z(_00385_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08378_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[26][17] ),
    .I1(_02337_),
    .S(_03877_),
    .Z(_03885_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08379_ (.I(_03885_),
    .Z(_00386_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08380_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[26][18] ),
    .I1(_02339_),
    .S(_03877_),
    .Z(_03886_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08381_ (.I(_03886_),
    .Z(_00387_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08382_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[26][19] ),
    .I1(_02341_),
    .S(_03877_),
    .Z(_03887_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08383_ (.I(_03887_),
    .Z(_00388_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08384_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[26][20] ),
    .I1(_02343_),
    .S(_03865_),
    .Z(_03888_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08385_ (.I(_03888_),
    .Z(_00389_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08386_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[26][21] ),
    .I1(_02260_),
    .S(_03865_),
    .Z(_03889_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08387_ (.I(_03889_),
    .Z(_00390_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08388_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[26][22] ),
    .I1(_02262_),
    .S(_03865_),
    .Z(_03890_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08389_ (.I(_03890_),
    .Z(_00391_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08390_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[26][23] ),
    .I1(_02264_),
    .S(_03865_),
    .Z(_03891_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08391_ (.I(_03891_),
    .Z(_00392_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08392_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[26][24] ),
    .I1(_02266_),
    .S(_03865_),
    .Z(_03892_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08393_ (.I(_03892_),
    .Z(_00393_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08394_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[26][25] ),
    .I1(_02268_),
    .S(_03865_),
    .Z(_03893_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08395_ (.I(_03893_),
    .Z(_00394_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08396_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[26][26] ),
    .I1(_02270_),
    .S(_03865_),
    .Z(_03894_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08397_ (.I(_03894_),
    .Z(_00395_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08398_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[26][27] ),
    .I1(_02351_),
    .S(_03865_),
    .Z(_03895_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08399_ (.I(_03895_),
    .Z(_00396_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08400_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[26][28] ),
    .I1(_02353_),
    .S(_03865_),
    .Z(_03896_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08401_ (.I(_03896_),
    .Z(_00397_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08402_ (.A1(_01441_),
    .A2(_03863_),
    .ZN(_03897_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _08403_ (.I(_03897_),
    .Z(_03898_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _08404_ (.I(_03898_),
    .Z(_03899_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08405_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[27][0] ),
    .I1(_02310_),
    .S(_03899_),
    .Z(_03900_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08406_ (.I(_03900_),
    .Z(_00398_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08407_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[27][1] ),
    .I1(_02393_),
    .S(_03899_),
    .Z(_03901_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08408_ (.I(_03901_),
    .Z(_00399_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08409_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[27][2] ),
    .I1(_02395_),
    .S(_03899_),
    .Z(_03902_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08410_ (.I(_03902_),
    .Z(_00400_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08411_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[27][3] ),
    .I1(_02397_),
    .S(_03899_),
    .Z(_03903_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08412_ (.I(_03903_),
    .Z(_00401_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08413_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[27][4] ),
    .I1(_02399_),
    .S(_03899_),
    .Z(_03904_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08414_ (.I(_03904_),
    .Z(_00402_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08415_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[27][5] ),
    .I1(_02401_),
    .S(_03899_),
    .Z(_03905_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08416_ (.I(_03905_),
    .Z(_00403_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08417_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[27][6] ),
    .I1(_02403_),
    .S(_03899_),
    .Z(_03906_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08418_ (.I(_03906_),
    .Z(_00404_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08419_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[27][7] ),
    .I1(_02405_),
    .S(_03899_),
    .Z(_03907_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08420_ (.I(_03907_),
    .Z(_00405_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08421_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[27][8] ),
    .I1(_02407_),
    .S(_03899_),
    .Z(_03908_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08422_ (.I(_03908_),
    .Z(_00406_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08423_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[27][9] ),
    .I1(_02409_),
    .S(_03899_),
    .Z(_03909_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08424_ (.I(_03909_),
    .Z(_00407_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _08425_ (.I(_03897_),
    .Z(_03910_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08426_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[27][10] ),
    .I1(_02411_),
    .S(_03910_),
    .Z(_03911_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08427_ (.I(_03911_),
    .Z(_00408_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08428_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[27][11] ),
    .I1(_02414_),
    .S(_03910_),
    .Z(_03912_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08429_ (.I(_03912_),
    .Z(_00409_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08430_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[27][12] ),
    .I1(_02242_),
    .S(_03910_),
    .Z(_03913_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08431_ (.I(_03913_),
    .Z(_00410_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08432_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[27][13] ),
    .I1(_02244_),
    .S(_03910_),
    .Z(_03914_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08433_ (.I(_03914_),
    .Z(_00411_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08434_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[27][14] ),
    .I1(_02246_),
    .S(_03910_),
    .Z(_03915_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08435_ (.I(_03915_),
    .Z(_00412_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08436_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[27][15] ),
    .I1(_02248_),
    .S(_03910_),
    .Z(_03916_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08437_ (.I(_03916_),
    .Z(_00413_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08438_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[27][16] ),
    .I1(_02335_),
    .S(_03910_),
    .Z(_03917_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08439_ (.I(_03917_),
    .Z(_00414_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08440_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[27][17] ),
    .I1(_02337_),
    .S(_03910_),
    .Z(_03918_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08441_ (.I(_03918_),
    .Z(_00415_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08442_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[27][18] ),
    .I1(_02339_),
    .S(_03910_),
    .Z(_03919_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08443_ (.I(_03919_),
    .Z(_00416_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08444_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[27][19] ),
    .I1(_02341_),
    .S(_03910_),
    .Z(_03920_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08445_ (.I(_03920_),
    .Z(_00417_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08446_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[27][20] ),
    .I1(_02343_),
    .S(_03898_),
    .Z(_03921_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08447_ (.I(_03921_),
    .Z(_00418_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08448_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[27][21] ),
    .I1(_02260_),
    .S(_03898_),
    .Z(_03922_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08449_ (.I(_03922_),
    .Z(_00419_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08450_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[27][22] ),
    .I1(_02262_),
    .S(_03898_),
    .Z(_03923_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08451_ (.I(_03923_),
    .Z(_00420_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08452_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[27][23] ),
    .I1(_02264_),
    .S(_03898_),
    .Z(_03924_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08453_ (.I(_03924_),
    .Z(_00421_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08454_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[27][24] ),
    .I1(_02266_),
    .S(_03898_),
    .Z(_03925_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08455_ (.I(_03925_),
    .Z(_00422_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08456_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[27][25] ),
    .I1(_02268_),
    .S(_03898_),
    .Z(_03926_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08457_ (.I(_03926_),
    .Z(_00423_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08458_ (.I(\soc.spi_video_ram_1.fifo_in_address[10] ),
    .Z(_03927_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08459_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[27][26] ),
    .I1(_03927_),
    .S(_03898_),
    .Z(_03928_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08460_ (.I(_03928_),
    .Z(_00424_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08461_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[27][27] ),
    .I1(_02351_),
    .S(_03898_),
    .Z(_03929_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08462_ (.I(_03929_),
    .Z(_00425_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08463_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[27][28] ),
    .I1(_02353_),
    .S(_03898_),
    .Z(_03930_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08464_ (.I(_03930_),
    .Z(_00426_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _08465_ (.A1(_02115_),
    .A2(_02312_),
    .A3(_03862_),
    .ZN(_03931_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08466_ (.A1(_03931_),
    .A2(_02214_),
    .ZN(_03932_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _08467_ (.I(_03932_),
    .Z(_03933_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _08468_ (.I(_03933_),
    .Z(_03934_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08469_ (.I0(_02113_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[28][0] ),
    .S(_03934_),
    .Z(_03935_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08470_ (.I(_03935_),
    .Z(_00427_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08471_ (.I0(_02122_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[28][1] ),
    .S(_03934_),
    .Z(_03936_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08472_ (.I(_03936_),
    .Z(_00428_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08473_ (.I0(_02124_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[28][2] ),
    .S(_03934_),
    .Z(_03937_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08474_ (.I(_03937_),
    .Z(_00429_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08475_ (.I0(_02126_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[28][3] ),
    .S(_03934_),
    .Z(_03938_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08476_ (.I(_03938_),
    .Z(_00430_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08477_ (.I0(_02128_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[28][4] ),
    .S(_03934_),
    .Z(_03939_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08478_ (.I(_03939_),
    .Z(_00431_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08479_ (.I0(_02130_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[28][5] ),
    .S(_03934_),
    .Z(_03940_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08480_ (.I(_03940_),
    .Z(_00432_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08481_ (.I0(_02132_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[28][6] ),
    .S(_03934_),
    .Z(_03941_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08482_ (.I(_03941_),
    .Z(_00433_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08483_ (.I0(_02134_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[28][7] ),
    .S(_03934_),
    .Z(_03942_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08484_ (.I(_03942_),
    .Z(_00434_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08485_ (.I0(_02136_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[28][8] ),
    .S(_03934_),
    .Z(_03943_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08486_ (.I(_03943_),
    .Z(_00435_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08487_ (.I0(_02138_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[28][9] ),
    .S(_03934_),
    .Z(_03944_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08488_ (.I(_03944_),
    .Z(_00436_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _08489_ (.I(_03932_),
    .Z(_03945_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08490_ (.I0(_02140_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[28][10] ),
    .S(_03945_),
    .Z(_03946_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08491_ (.I(_03946_),
    .Z(_00437_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08492_ (.I0(_02143_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[28][11] ),
    .S(_03945_),
    .Z(_03947_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08493_ (.I(_03947_),
    .Z(_00438_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08494_ (.I0(_02145_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[28][12] ),
    .S(_03945_),
    .Z(_03948_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08495_ (.I(_03948_),
    .Z(_00439_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08496_ (.I0(_02147_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[28][13] ),
    .S(_03945_),
    .Z(_03949_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08497_ (.I(_03949_),
    .Z(_00440_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08498_ (.I0(_02149_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[28][14] ),
    .S(_03945_),
    .Z(_03950_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08499_ (.I(_03950_),
    .Z(_00441_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08500_ (.I0(_02151_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[28][15] ),
    .S(_03945_),
    .Z(_03951_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08501_ (.I(_03951_),
    .Z(_00442_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08502_ (.I0(_02153_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[28][16] ),
    .S(_03945_),
    .Z(_03952_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08503_ (.I(_03952_),
    .Z(_00443_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08504_ (.I0(_02155_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[28][17] ),
    .S(_03945_),
    .Z(_03953_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08505_ (.I(_03953_),
    .Z(_00444_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08506_ (.I0(_02157_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[28][18] ),
    .S(_03945_),
    .Z(_03954_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08507_ (.I(_03954_),
    .Z(_00445_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08508_ (.I0(_02159_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[28][19] ),
    .S(_03945_),
    .Z(_03955_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08509_ (.I(_03955_),
    .Z(_00446_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08510_ (.I0(_02161_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[28][20] ),
    .S(_03933_),
    .Z(_03956_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08511_ (.I(_03956_),
    .Z(_00447_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08512_ (.I0(_02163_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[28][21] ),
    .S(_03933_),
    .Z(_03957_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08513_ (.I(_03957_),
    .Z(_00448_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08514_ (.I0(_02165_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[28][22] ),
    .S(_03933_),
    .Z(_03958_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08515_ (.I(_03958_),
    .Z(_00449_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08516_ (.I0(_02167_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[28][23] ),
    .S(_03933_),
    .Z(_03959_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08517_ (.I(_03959_),
    .Z(_00450_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08518_ (.I0(_02169_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[28][24] ),
    .S(_03933_),
    .Z(_03960_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08519_ (.I(_03960_),
    .Z(_00451_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08520_ (.I0(_02171_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[28][25] ),
    .S(_03933_),
    .Z(_03961_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08521_ (.I(_03961_),
    .Z(_00452_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08522_ (.I0(_02173_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[28][26] ),
    .S(_03933_),
    .Z(_03962_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08523_ (.I(_03962_),
    .Z(_00453_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08524_ (.I0(_02175_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[28][27] ),
    .S(_03933_),
    .Z(_03963_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08525_ (.I(_03963_),
    .Z(_00454_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08526_ (.I0(_02177_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[28][28] ),
    .S(_03933_),
    .Z(_03964_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08527_ (.I(_03964_),
    .Z(_00455_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08528_ (.A1(_02114_),
    .A2(_02276_),
    .ZN(_03965_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _08529_ (.I(_03965_),
    .Z(_03966_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _08530_ (.I(_03966_),
    .Z(_03967_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08531_ (.I0(_02113_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[2][0] ),
    .S(_03967_),
    .Z(_03968_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08532_ (.I(_03968_),
    .Z(_00456_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08533_ (.I0(_02122_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[2][1] ),
    .S(_03967_),
    .Z(_03969_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08534_ (.I(_03969_),
    .Z(_00457_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08535_ (.I0(_02124_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[2][2] ),
    .S(_03967_),
    .Z(_03970_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08536_ (.I(_03970_),
    .Z(_00458_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08537_ (.I0(_02126_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[2][3] ),
    .S(_03967_),
    .Z(_03971_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08538_ (.I(_03971_),
    .Z(_00459_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08539_ (.I0(_02128_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[2][4] ),
    .S(_03967_),
    .Z(_03972_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08540_ (.I(_03972_),
    .Z(_00460_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08541_ (.I0(_02130_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[2][5] ),
    .S(_03967_),
    .Z(_03973_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08542_ (.I(_03973_),
    .Z(_00461_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08543_ (.I0(_02132_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[2][6] ),
    .S(_03967_),
    .Z(_03974_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08544_ (.I(_03974_),
    .Z(_00462_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08545_ (.I0(_02134_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[2][7] ),
    .S(_03967_),
    .Z(_03975_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08546_ (.I(_03975_),
    .Z(_00463_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08547_ (.I0(_02136_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[2][8] ),
    .S(_03967_),
    .Z(_03976_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08548_ (.I(_03976_),
    .Z(_00464_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08549_ (.I0(_02138_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[2][9] ),
    .S(_03967_),
    .Z(_03977_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08550_ (.I(_03977_),
    .Z(_00465_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _08551_ (.I(_03965_),
    .Z(_03978_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08552_ (.I0(_02140_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[2][10] ),
    .S(_03978_),
    .Z(_03979_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08553_ (.I(_03979_),
    .Z(_00466_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08554_ (.I0(_02143_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[2][11] ),
    .S(_03978_),
    .Z(_03980_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08555_ (.I(_03980_),
    .Z(_00467_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08556_ (.I0(_02145_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[2][12] ),
    .S(_03978_),
    .Z(_03981_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08557_ (.I(_03981_),
    .Z(_00468_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08558_ (.I0(_02147_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[2][13] ),
    .S(_03978_),
    .Z(_03982_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08559_ (.I(_03982_),
    .Z(_00469_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08560_ (.I0(_02149_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[2][14] ),
    .S(_03978_),
    .Z(_03983_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08561_ (.I(_03983_),
    .Z(_00470_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08562_ (.I0(_02151_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[2][15] ),
    .S(_03978_),
    .Z(_03984_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08563_ (.I(_03984_),
    .Z(_00471_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08564_ (.I0(_02153_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[2][16] ),
    .S(_03978_),
    .Z(_03985_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08565_ (.I(_03985_),
    .Z(_00472_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08566_ (.I0(_02155_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[2][17] ),
    .S(_03978_),
    .Z(_03986_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08567_ (.I(_03986_),
    .Z(_00473_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08568_ (.I0(_02157_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[2][18] ),
    .S(_03978_),
    .Z(_03987_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08569_ (.I(_03987_),
    .Z(_00474_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08570_ (.I0(_02159_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[2][19] ),
    .S(_03978_),
    .Z(_03988_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08571_ (.I(_03988_),
    .Z(_00475_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08572_ (.I0(_02161_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[2][20] ),
    .S(_03966_),
    .Z(_03989_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08573_ (.I(_03989_),
    .Z(_00476_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08574_ (.I0(_02163_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[2][21] ),
    .S(_03966_),
    .Z(_03990_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08575_ (.I(_03990_),
    .Z(_00477_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08576_ (.I0(_02165_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[2][22] ),
    .S(_03966_),
    .Z(_03991_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08577_ (.I(_03991_),
    .Z(_00478_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08578_ (.I0(_02167_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[2][23] ),
    .S(_03966_),
    .Z(_03992_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08579_ (.I(_03992_),
    .Z(_00479_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08580_ (.I0(_02169_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[2][24] ),
    .S(_03966_),
    .Z(_03993_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08581_ (.I(_03993_),
    .Z(_00480_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08582_ (.I0(_02171_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[2][25] ),
    .S(_03966_),
    .Z(_03994_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08583_ (.I(_03994_),
    .Z(_00481_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08584_ (.I0(_02173_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[2][26] ),
    .S(_03966_),
    .Z(_03995_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08585_ (.I(_03995_),
    .Z(_00482_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08586_ (.I0(_02175_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[2][27] ),
    .S(_03966_),
    .Z(_03996_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08587_ (.I(_03996_),
    .Z(_00483_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08588_ (.I0(_02177_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[2][28] ),
    .S(_03966_),
    .Z(_03997_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08589_ (.I(_03997_),
    .Z(_00484_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08590_ (.A1(_03931_),
    .A2(_02114_),
    .ZN(_03998_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _08591_ (.I(_03998_),
    .Z(_03999_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _08592_ (.I(_03999_),
    .Z(_04000_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08593_ (.I0(_02113_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[30][0] ),
    .S(_04000_),
    .Z(_04001_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08594_ (.I(_04001_),
    .Z(_00485_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08595_ (.I0(_02122_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[30][1] ),
    .S(_04000_),
    .Z(_04002_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08596_ (.I(_04002_),
    .Z(_00486_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08597_ (.I0(_02124_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[30][2] ),
    .S(_04000_),
    .Z(_04003_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08598_ (.I(_04003_),
    .Z(_00487_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08599_ (.I0(_02126_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[30][3] ),
    .S(_04000_),
    .Z(_04004_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08600_ (.I(_04004_),
    .Z(_00488_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08601_ (.I0(_02128_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[30][4] ),
    .S(_04000_),
    .Z(_04005_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08602_ (.I(_04005_),
    .Z(_00489_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08603_ (.I0(_02130_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[30][5] ),
    .S(_04000_),
    .Z(_04006_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08604_ (.I(_04006_),
    .Z(_00490_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08605_ (.I0(_02132_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[30][6] ),
    .S(_04000_),
    .Z(_04007_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08606_ (.I(_04007_),
    .Z(_00491_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08607_ (.I0(_02134_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[30][7] ),
    .S(_04000_),
    .Z(_04008_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08608_ (.I(_04008_),
    .Z(_00492_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08609_ (.I0(_02136_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[30][8] ),
    .S(_04000_),
    .Z(_04009_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08610_ (.I(_04009_),
    .Z(_00493_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08611_ (.I0(_02138_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[30][9] ),
    .S(_04000_),
    .Z(_04010_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08612_ (.I(_04010_),
    .Z(_00494_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _08613_ (.I(_03998_),
    .Z(_04011_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08614_ (.I0(_02140_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[30][10] ),
    .S(_04011_),
    .Z(_04012_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08615_ (.I(_04012_),
    .Z(_00495_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08616_ (.I0(_02143_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[30][11] ),
    .S(_04011_),
    .Z(_04013_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08617_ (.I(_04013_),
    .Z(_00496_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08618_ (.I0(_02145_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[30][12] ),
    .S(_04011_),
    .Z(_04014_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08619_ (.I(_04014_),
    .Z(_00497_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08620_ (.I0(_02147_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[30][13] ),
    .S(_04011_),
    .Z(_04015_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08621_ (.I(_04015_),
    .Z(_00498_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08622_ (.I0(_02149_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[30][14] ),
    .S(_04011_),
    .Z(_04016_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08623_ (.I(_04016_),
    .Z(_00499_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08624_ (.I0(_02151_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[30][15] ),
    .S(_04011_),
    .Z(_04017_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08625_ (.I(_04017_),
    .Z(_00500_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08626_ (.I0(_02153_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[30][16] ),
    .S(_04011_),
    .Z(_04018_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08627_ (.I(_04018_),
    .Z(_00501_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08628_ (.I0(_02155_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[30][17] ),
    .S(_04011_),
    .Z(_04019_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08629_ (.I(_04019_),
    .Z(_00502_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08630_ (.I0(_02157_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[30][18] ),
    .S(_04011_),
    .Z(_04020_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08631_ (.I(_04020_),
    .Z(_00503_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08632_ (.I0(_02159_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[30][19] ),
    .S(_04011_),
    .Z(_04021_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08633_ (.I(_04021_),
    .Z(_00504_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08634_ (.I0(_02161_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[30][20] ),
    .S(_03999_),
    .Z(_04022_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08635_ (.I(_04022_),
    .Z(_00505_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08636_ (.I0(_02163_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[30][21] ),
    .S(_03999_),
    .Z(_04023_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08637_ (.I(_04023_),
    .Z(_00506_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08638_ (.I0(_02165_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[30][22] ),
    .S(_03999_),
    .Z(_04024_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08639_ (.I(_04024_),
    .Z(_00507_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08640_ (.I0(_02167_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[30][23] ),
    .S(_03999_),
    .Z(_04025_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08641_ (.I(_04025_),
    .Z(_00508_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08642_ (.I0(_02169_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[30][24] ),
    .S(_03999_),
    .Z(_04026_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08643_ (.I(_04026_),
    .Z(_00509_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08644_ (.I0(_02171_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[30][25] ),
    .S(_03999_),
    .Z(_04027_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08645_ (.I(_04027_),
    .Z(_00510_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08646_ (.I0(_02173_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[30][26] ),
    .S(_03999_),
    .Z(_04028_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08647_ (.I(_04028_),
    .Z(_00511_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08648_ (.I0(_02175_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[30][27] ),
    .S(_03999_),
    .Z(_04029_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08649_ (.I(_04029_),
    .Z(_00512_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08650_ (.I0(_02177_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[30][28] ),
    .S(_03999_),
    .Z(_04030_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08651_ (.I(_04030_),
    .Z(_00513_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _08652_ (.A1(\soc.spi_video_ram_1.write_fifo.write_pointer[4] ),
    .A2(_01449_),
    .ZN(_04031_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _08653_ (.I(_04031_),
    .Z(_04032_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08654_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[15][0] ),
    .I1(_02310_),
    .S(_04032_),
    .Z(_04033_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08655_ (.I(_04033_),
    .Z(_00514_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08656_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[15][1] ),
    .I1(_02393_),
    .S(_04032_),
    .Z(_04034_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08657_ (.I(_04034_),
    .Z(_00515_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08658_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[15][2] ),
    .I1(_02395_),
    .S(_04032_),
    .Z(_04035_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08659_ (.I(_04035_),
    .Z(_00516_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08660_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[15][3] ),
    .I1(_02397_),
    .S(_04032_),
    .Z(_04036_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08661_ (.I(_04036_),
    .Z(_00517_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08662_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[15][4] ),
    .I1(_02399_),
    .S(_04032_),
    .Z(_04037_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08663_ (.I(_04037_),
    .Z(_00518_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08664_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[15][5] ),
    .I1(_02401_),
    .S(_04032_),
    .Z(_04038_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08665_ (.I(_04038_),
    .Z(_00519_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08666_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[15][6] ),
    .I1(_02403_),
    .S(_04032_),
    .Z(_04039_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08667_ (.I(_04039_),
    .Z(_00520_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08668_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[15][7] ),
    .I1(_02405_),
    .S(_04032_),
    .Z(_04040_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08669_ (.I(_04040_),
    .Z(_00521_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08670_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[15][8] ),
    .I1(_02407_),
    .S(_04032_),
    .Z(_04041_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08671_ (.I(_04041_),
    .Z(_00522_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08672_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[15][9] ),
    .I1(_02409_),
    .S(_04032_),
    .Z(_04042_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08673_ (.I(_04042_),
    .Z(_00523_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _08674_ (.I(_04031_),
    .Z(_04043_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08675_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[15][10] ),
    .I1(_02411_),
    .S(_04043_),
    .Z(_04044_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08676_ (.I(_04044_),
    .Z(_00524_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08677_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[15][11] ),
    .I1(_02414_),
    .S(_04043_),
    .Z(_04045_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08678_ (.I(_04045_),
    .Z(_00525_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08679_ (.I(_04043_),
    .Z(_04046_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08680_ (.I(\soc.spi_video_ram_1.fifo_in_data[12] ),
    .Z(_04047_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08681_ (.I(_04031_),
    .Z(_04048_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08682_ (.A1(_04047_),
    .A2(_04048_),
    .ZN(_04049_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08683_ (.A1(_03140_),
    .A2(_04046_),
    .B(_04049_),
    .ZN(_00526_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08684_ (.I(\soc.spi_video_ram_1.fifo_in_data[13] ),
    .Z(_04050_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08685_ (.A1(_04050_),
    .A2(_04048_),
    .ZN(_04051_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08686_ (.A1(_03214_),
    .A2(_04046_),
    .B(_04051_),
    .ZN(_00527_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08687_ (.I(\soc.spi_video_ram_1.fifo_in_data[14] ),
    .Z(_04052_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08688_ (.A1(_04052_),
    .A2(_04048_),
    .ZN(_04053_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08689_ (.A1(_03312_),
    .A2(_04046_),
    .B(_04053_),
    .ZN(_00528_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08690_ (.I(\soc.spi_video_ram_1.fifo_in_data[15] ),
    .Z(_04054_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08691_ (.A1(_04054_),
    .A2(_04048_),
    .ZN(_04055_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08692_ (.A1(_03404_),
    .A2(_04046_),
    .B(_04055_),
    .ZN(_00529_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08693_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[15][16] ),
    .I1(_02335_),
    .S(_04043_),
    .Z(_04056_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08694_ (.I(_04056_),
    .Z(_00530_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08695_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[15][17] ),
    .I1(_02337_),
    .S(_04043_),
    .Z(_04057_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08696_ (.I(_04057_),
    .Z(_00531_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08697_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[15][18] ),
    .I1(_02339_),
    .S(_04043_),
    .Z(_04058_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08698_ (.I(_04058_),
    .Z(_00532_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08699_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[15][19] ),
    .I1(_02341_),
    .S(_04043_),
    .Z(_04059_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08700_ (.I(_04059_),
    .Z(_00533_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08701_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[15][20] ),
    .I1(_02343_),
    .S(_04043_),
    .Z(_04060_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08702_ (.I(_04060_),
    .Z(_00534_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08703_ (.I(\soc.spi_video_ram_1.fifo_in_address[5] ),
    .Z(_04061_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08704_ (.A1(_04061_),
    .A2(_04048_),
    .ZN(_04062_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08705_ (.A1(_03541_),
    .A2(_04046_),
    .B(_04062_),
    .ZN(_00535_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08706_ (.I(\soc.spi_video_ram_1.fifo_in_address[6] ),
    .Z(_04063_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08707_ (.A1(_04063_),
    .A2(_04048_),
    .ZN(_04064_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08708_ (.A1(_03511_),
    .A2(_04046_),
    .B(_04064_),
    .ZN(_00536_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08709_ (.I(\soc.spi_video_ram_1.fifo_in_address[7] ),
    .Z(_04065_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08710_ (.A1(_04065_),
    .A2(_04048_),
    .ZN(_04066_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08711_ (.A1(_03464_),
    .A2(_04046_),
    .B(_04066_),
    .ZN(_00537_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08712_ (.I(\soc.spi_video_ram_1.fifo_in_address[8] ),
    .Z(_04067_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08713_ (.A1(_04067_),
    .A2(_04048_),
    .ZN(_04068_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08714_ (.A1(_03368_),
    .A2(_04046_),
    .B(_04068_),
    .ZN(_00538_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08715_ (.I(\soc.spi_video_ram_1.fifo_in_address[9] ),
    .Z(_04069_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08716_ (.A1(_04069_),
    .A2(_04048_),
    .ZN(_04070_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08717_ (.A1(_03270_),
    .A2(_04046_),
    .B(_04070_),
    .ZN(_00539_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08718_ (.A1(_03927_),
    .A2(_04048_),
    .ZN(_04071_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08719_ (.A1(_03169_),
    .A2(_04046_),
    .B(_04071_),
    .ZN(_00540_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08720_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[15][27] ),
    .I1(_02351_),
    .S(_04043_),
    .Z(_04072_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08721_ (.I(_04072_),
    .Z(_00541_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08722_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[15][28] ),
    .I1(_02353_),
    .S(_04043_),
    .Z(_04073_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08723_ (.I(_04073_),
    .Z(_00542_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _08724_ (.A1(\soc.spi_video_ram_1.write_fifo.write_pointer[1] ),
    .A2(_01405_),
    .A3(_03863_),
    .ZN(_04074_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _08725_ (.I(_04074_),
    .Z(_04075_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _08726_ (.I(_04075_),
    .Z(_04076_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08727_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[24][0] ),
    .I1(_02310_),
    .S(_04076_),
    .Z(_04077_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08728_ (.I(_04077_),
    .Z(_00543_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08729_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[24][1] ),
    .I1(_02393_),
    .S(_04076_),
    .Z(_04078_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08730_ (.I(_04078_),
    .Z(_00544_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08731_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[24][2] ),
    .I1(_02395_),
    .S(_04076_),
    .Z(_04079_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08732_ (.I(_04079_),
    .Z(_00545_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08733_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[24][3] ),
    .I1(_02397_),
    .S(_04076_),
    .Z(_04080_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08734_ (.I(_04080_),
    .Z(_00546_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08735_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[24][4] ),
    .I1(_02399_),
    .S(_04076_),
    .Z(_04081_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08736_ (.I(_04081_),
    .Z(_00547_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08737_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[24][5] ),
    .I1(_02401_),
    .S(_04076_),
    .Z(_04082_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08738_ (.I(_04082_),
    .Z(_00548_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08739_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[24][6] ),
    .I1(_02403_),
    .S(_04076_),
    .Z(_04083_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08740_ (.I(_04083_),
    .Z(_00549_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08741_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[24][7] ),
    .I1(_02405_),
    .S(_04076_),
    .Z(_04084_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08742_ (.I(_04084_),
    .Z(_00550_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08743_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[24][8] ),
    .I1(_02407_),
    .S(_04076_),
    .Z(_04085_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08744_ (.I(_04085_),
    .Z(_00551_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08745_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[24][9] ),
    .I1(_02409_),
    .S(_04076_),
    .Z(_04086_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08746_ (.I(_04086_),
    .Z(_00552_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _08747_ (.I(_04074_),
    .Z(_04087_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08748_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[24][10] ),
    .I1(_02411_),
    .S(_04087_),
    .Z(_04088_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08749_ (.I(_04088_),
    .Z(_00553_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08750_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[24][11] ),
    .I1(_02414_),
    .S(_04087_),
    .Z(_04089_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08751_ (.I(_04089_),
    .Z(_00554_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08752_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[24][12] ),
    .I1(_04047_),
    .S(_04087_),
    .Z(_04090_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08753_ (.I(_04090_),
    .Z(_00555_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08754_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[24][13] ),
    .I1(_04050_),
    .S(_04087_),
    .Z(_04091_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08755_ (.I(_04091_),
    .Z(_00556_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08756_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[24][14] ),
    .I1(_04052_),
    .S(_04087_),
    .Z(_04092_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08757_ (.I(_04092_),
    .Z(_00557_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08758_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[24][15] ),
    .I1(_04054_),
    .S(_04087_),
    .Z(_04093_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08759_ (.I(_04093_),
    .Z(_00558_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08760_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[24][16] ),
    .I1(_02335_),
    .S(_04087_),
    .Z(_04094_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08761_ (.I(_04094_),
    .Z(_00559_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08762_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[24][17] ),
    .I1(_02337_),
    .S(_04087_),
    .Z(_04095_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08763_ (.I(_04095_),
    .Z(_00560_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08764_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[24][18] ),
    .I1(_02339_),
    .S(_04087_),
    .Z(_04096_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08765_ (.I(_04096_),
    .Z(_00561_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08766_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[24][19] ),
    .I1(_02341_),
    .S(_04087_),
    .Z(_04097_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08767_ (.I(_04097_),
    .Z(_00562_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08768_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[24][20] ),
    .I1(_02343_),
    .S(_04075_),
    .Z(_04098_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08769_ (.I(_04098_),
    .Z(_00563_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08770_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[24][21] ),
    .I1(_04061_),
    .S(_04075_),
    .Z(_04099_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08771_ (.I(_04099_),
    .Z(_00564_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08772_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[24][22] ),
    .I1(_04063_),
    .S(_04075_),
    .Z(_04100_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08773_ (.I(_04100_),
    .Z(_00565_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08774_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[24][23] ),
    .I1(_04065_),
    .S(_04075_),
    .Z(_04101_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08775_ (.I(_04101_),
    .Z(_00566_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08776_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[24][24] ),
    .I1(_04067_),
    .S(_04075_),
    .Z(_04102_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08777_ (.I(_04102_),
    .Z(_00567_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08778_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[24][25] ),
    .I1(_04069_),
    .S(_04075_),
    .Z(_04103_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08779_ (.I(_04103_),
    .Z(_00568_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08780_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[24][26] ),
    .I1(_03927_),
    .S(_04075_),
    .Z(_04104_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08781_ (.I(_04104_),
    .Z(_00569_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08782_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[24][27] ),
    .I1(_02351_),
    .S(_04075_),
    .Z(_04105_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08783_ (.I(_04105_),
    .Z(_00570_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08784_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[24][28] ),
    .I1(_02353_),
    .S(_04075_),
    .Z(_04106_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08785_ (.I(_04106_),
    .Z(_00571_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08786_ (.A1(_02115_),
    .A2(_01403_),
    .ZN(_04107_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08787_ (.A1(_02116_),
    .A2(_01445_),
    .A3(_04107_),
    .ZN(_04108_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _08788_ (.I(_04108_),
    .Z(_04109_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _08789_ (.I(_04109_),
    .Z(_04110_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08790_ (.I0(_02113_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[23][0] ),
    .S(_04110_),
    .Z(_04111_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08791_ (.I(_04111_),
    .Z(_00572_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08792_ (.I0(_02122_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[23][1] ),
    .S(_04110_),
    .Z(_04112_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08793_ (.I(_04112_),
    .Z(_00573_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08794_ (.I0(_02124_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[23][2] ),
    .S(_04110_),
    .Z(_04113_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08795_ (.I(_04113_),
    .Z(_00574_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08796_ (.I0(_02126_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[23][3] ),
    .S(_04110_),
    .Z(_04114_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08797_ (.I(_04114_),
    .Z(_00575_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08798_ (.I0(_02128_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[23][4] ),
    .S(_04110_),
    .Z(_04115_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08799_ (.I(_04115_),
    .Z(_00576_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08800_ (.I0(_02130_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[23][5] ),
    .S(_04110_),
    .Z(_04116_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08801_ (.I(_04116_),
    .Z(_00577_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _08802_ (.I(_04109_),
    .Z(_04117_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08803_ (.I0(_02132_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[23][6] ),
    .S(_04117_),
    .Z(_04118_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08804_ (.I(_04118_),
    .Z(_00578_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08805_ (.I0(_02134_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[23][7] ),
    .S(_04117_),
    .Z(_04119_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08806_ (.I(_04119_),
    .Z(_00579_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08807_ (.I0(_02136_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[23][8] ),
    .S(_04117_),
    .Z(_04120_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08808_ (.I(_04120_),
    .Z(_00580_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08809_ (.I0(_02138_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[23][9] ),
    .S(_04117_),
    .Z(_04121_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08810_ (.I(_04121_),
    .Z(_00581_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08811_ (.I0(_02140_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[23][10] ),
    .S(_04117_),
    .Z(_04122_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08812_ (.I(_04122_),
    .Z(_00582_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08813_ (.I0(_02143_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[23][11] ),
    .S(_04117_),
    .Z(_04123_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08814_ (.I(_04123_),
    .Z(_00583_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08815_ (.I(_04109_),
    .Z(_04124_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08816_ (.A1(_04047_),
    .A2(_04124_),
    .ZN(_04125_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08817_ (.A1(_03109_),
    .A2(_04124_),
    .B(_04125_),
    .ZN(_00584_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08818_ (.I0(_02147_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[23][13] ),
    .S(_04117_),
    .Z(_04126_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08819_ (.I(_04126_),
    .Z(_00585_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08820_ (.I0(_02149_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[23][14] ),
    .S(_04117_),
    .Z(_04127_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08821_ (.I(_04127_),
    .Z(_00586_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08822_ (.I0(_02151_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[23][15] ),
    .S(_04117_),
    .Z(_04128_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08823_ (.I(_04128_),
    .Z(_00587_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08824_ (.I0(_02153_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[23][16] ),
    .S(_04117_),
    .Z(_04129_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08825_ (.I(_04129_),
    .Z(_00588_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08826_ (.I0(_02155_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[23][17] ),
    .S(_04109_),
    .Z(_04130_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08827_ (.I(_04130_),
    .Z(_00589_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08828_ (.I0(_02157_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[23][18] ),
    .S(_04109_),
    .Z(_04131_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08829_ (.I(_04131_),
    .Z(_00590_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08830_ (.I0(_02159_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[23][19] ),
    .S(_04109_),
    .Z(_04132_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08831_ (.I(_04132_),
    .Z(_00591_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08832_ (.I0(_02161_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[23][20] ),
    .S(_04109_),
    .Z(_04133_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08833_ (.I(_04133_),
    .Z(_00592_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08834_ (.A1(_04061_),
    .A2(_04124_),
    .ZN(_04134_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08835_ (.A1(_03554_),
    .A2(_04124_),
    .B(_04134_),
    .ZN(_00593_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08836_ (.A1(_04063_),
    .A2(_04124_),
    .ZN(_04135_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08837_ (.A1(_03482_),
    .A2(_04124_),
    .B(_04135_),
    .ZN(_00594_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08838_ (.A1(_04065_),
    .A2(_04110_),
    .ZN(_04136_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08839_ (.A1(_03431_),
    .A2(_04124_),
    .B(_04136_),
    .ZN(_00595_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08840_ (.A1(_04067_),
    .A2(_04110_),
    .ZN(_04137_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08841_ (.A1(_03335_),
    .A2(_04124_),
    .B(_04137_),
    .ZN(_00596_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08842_ (.A1(_04069_),
    .A2(_04110_),
    .ZN(_04138_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08843_ (.A1(_03237_),
    .A2(_04124_),
    .B(_04138_),
    .ZN(_00597_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08844_ (.A1(_03927_),
    .A2(_04110_),
    .ZN(_04139_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08845_ (.A1(_03151_),
    .A2(_04124_),
    .B(_04139_),
    .ZN(_00598_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08846_ (.I0(_02175_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[23][27] ),
    .S(_04109_),
    .Z(_04140_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08847_ (.I(_04140_),
    .Z(_00599_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08848_ (.I0(_02177_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[23][28] ),
    .S(_04109_),
    .Z(_04141_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08849_ (.I(_04141_),
    .Z(_00600_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08850_ (.A1(_02311_),
    .A2(_03863_),
    .ZN(_04142_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _08851_ (.I(_04142_),
    .Z(_04143_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _08852_ (.I(_04143_),
    .Z(_04144_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08853_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[25][0] ),
    .I1(_02310_),
    .S(_04144_),
    .Z(_04145_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08854_ (.I(_04145_),
    .Z(_00601_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08855_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[25][1] ),
    .I1(_02393_),
    .S(_04144_),
    .Z(_04146_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08856_ (.I(_04146_),
    .Z(_00602_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08857_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[25][2] ),
    .I1(_02395_),
    .S(_04144_),
    .Z(_04147_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08858_ (.I(_04147_),
    .Z(_00603_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08859_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[25][3] ),
    .I1(_02397_),
    .S(_04144_),
    .Z(_04148_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08860_ (.I(_04148_),
    .Z(_00604_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08861_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[25][4] ),
    .I1(_02399_),
    .S(_04144_),
    .Z(_04149_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08862_ (.I(_04149_),
    .Z(_00605_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08863_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[25][5] ),
    .I1(_02401_),
    .S(_04144_),
    .Z(_04150_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08864_ (.I(_04150_),
    .Z(_00606_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08865_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[25][6] ),
    .I1(_02403_),
    .S(_04144_),
    .Z(_04151_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08866_ (.I(_04151_),
    .Z(_00607_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08867_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[25][7] ),
    .I1(_02405_),
    .S(_04144_),
    .Z(_04152_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08868_ (.I(_04152_),
    .Z(_00608_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08869_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[25][8] ),
    .I1(_02407_),
    .S(_04144_),
    .Z(_04153_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08870_ (.I(_04153_),
    .Z(_00609_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08871_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[25][9] ),
    .I1(_02409_),
    .S(_04144_),
    .Z(_04154_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08872_ (.I(_04154_),
    .Z(_00610_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _08873_ (.I(_04142_),
    .Z(_04155_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08874_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[25][10] ),
    .I1(_02411_),
    .S(_04155_),
    .Z(_04156_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08875_ (.I(_04156_),
    .Z(_00611_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08876_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[25][11] ),
    .I1(_02414_),
    .S(_04155_),
    .Z(_04157_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08877_ (.I(_04157_),
    .Z(_00612_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08878_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[25][12] ),
    .I1(_04047_),
    .S(_04155_),
    .Z(_04158_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08879_ (.I(_04158_),
    .Z(_00613_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08880_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[25][13] ),
    .I1(_04050_),
    .S(_04155_),
    .Z(_04159_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08881_ (.I(_04159_),
    .Z(_00614_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08882_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[25][14] ),
    .I1(_04052_),
    .S(_04155_),
    .Z(_04160_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08883_ (.I(_04160_),
    .Z(_00615_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08884_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[25][15] ),
    .I1(_04054_),
    .S(_04155_),
    .Z(_04161_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08885_ (.I(_04161_),
    .Z(_00616_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08886_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[25][16] ),
    .I1(_02335_),
    .S(_04155_),
    .Z(_04162_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08887_ (.I(_04162_),
    .Z(_00617_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08888_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[25][17] ),
    .I1(_02337_),
    .S(_04155_),
    .Z(_04163_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08889_ (.I(_04163_),
    .Z(_00618_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08890_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[25][18] ),
    .I1(_02339_),
    .S(_04155_),
    .Z(_04164_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08891_ (.I(_04164_),
    .Z(_00619_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08892_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[25][19] ),
    .I1(_02341_),
    .S(_04155_),
    .Z(_04165_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08893_ (.I(_04165_),
    .Z(_00620_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08894_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[25][20] ),
    .I1(_02343_),
    .S(_04143_),
    .Z(_04166_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08895_ (.I(_04166_),
    .Z(_00621_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08896_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[25][21] ),
    .I1(_04061_),
    .S(_04143_),
    .Z(_04167_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08897_ (.I(_04167_),
    .Z(_00622_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08898_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[25][22] ),
    .I1(_04063_),
    .S(_04143_),
    .Z(_04168_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08899_ (.I(_04168_),
    .Z(_00623_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08900_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[25][23] ),
    .I1(_04065_),
    .S(_04143_),
    .Z(_04169_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08901_ (.I(_04169_),
    .Z(_00624_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08902_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[25][24] ),
    .I1(_04067_),
    .S(_04143_),
    .Z(_04170_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08903_ (.I(_04170_),
    .Z(_00625_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08904_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[25][25] ),
    .I1(_04069_),
    .S(_04143_),
    .Z(_04171_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08905_ (.I(_04171_),
    .Z(_00626_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08906_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[25][26] ),
    .I1(_03927_),
    .S(_04143_),
    .Z(_04172_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08907_ (.I(_04172_),
    .Z(_00627_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08908_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[25][27] ),
    .I1(_02351_),
    .S(_04143_),
    .Z(_04173_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08909_ (.I(_04173_),
    .Z(_00628_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08910_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[25][28] ),
    .I1(_02353_),
    .S(_04143_),
    .Z(_04174_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08911_ (.I(_04174_),
    .Z(_00629_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08912_ (.A1(_02116_),
    .A2(_04107_),
    .ZN(_04175_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08913_ (.A1(_02388_),
    .A2(_04175_),
    .ZN(_04176_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _08914_ (.I(_04176_),
    .Z(_04177_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _08915_ (.I(_04177_),
    .Z(_04178_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08916_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[22][0] ),
    .I1(_02310_),
    .S(_04178_),
    .Z(_04179_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08917_ (.I(_04179_),
    .Z(_00630_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08918_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[22][1] ),
    .I1(_02393_),
    .S(_04178_),
    .Z(_04180_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08919_ (.I(_04180_),
    .Z(_00631_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08920_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[22][2] ),
    .I1(_02395_),
    .S(_04178_),
    .Z(_04181_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08921_ (.I(_04181_),
    .Z(_00632_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08922_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[22][3] ),
    .I1(_02397_),
    .S(_04178_),
    .Z(_04182_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08923_ (.I(_04182_),
    .Z(_00633_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08924_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[22][4] ),
    .I1(_02399_),
    .S(_04178_),
    .Z(_04183_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08925_ (.I(_04183_),
    .Z(_00634_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08926_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[22][5] ),
    .I1(_02401_),
    .S(_04178_),
    .Z(_04184_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08927_ (.I(_04184_),
    .Z(_00635_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08928_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[22][6] ),
    .I1(_02403_),
    .S(_04178_),
    .Z(_04185_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08929_ (.I(_04185_),
    .Z(_00636_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08930_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[22][7] ),
    .I1(_02405_),
    .S(_04178_),
    .Z(_04186_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08931_ (.I(_04186_),
    .Z(_00637_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08932_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[22][8] ),
    .I1(_02407_),
    .S(_04178_),
    .Z(_04187_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08933_ (.I(_04187_),
    .Z(_00638_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08934_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[22][9] ),
    .I1(_02409_),
    .S(_04178_),
    .Z(_04188_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08935_ (.I(_04188_),
    .Z(_00639_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _08936_ (.I(_04176_),
    .Z(_04189_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08937_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[22][10] ),
    .I1(_02411_),
    .S(_04189_),
    .Z(_04190_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08938_ (.I(_04190_),
    .Z(_00640_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08939_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[22][11] ),
    .I1(_02414_),
    .S(_04189_),
    .Z(_04191_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08940_ (.I(_04191_),
    .Z(_00641_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08941_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[22][12] ),
    .I1(_04047_),
    .S(_04189_),
    .Z(_04192_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08942_ (.I(_04192_),
    .Z(_00642_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08943_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[22][13] ),
    .I1(_04050_),
    .S(_04189_),
    .Z(_04193_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08944_ (.I(_04193_),
    .Z(_00643_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08945_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[22][14] ),
    .I1(_04052_),
    .S(_04189_),
    .Z(_04194_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08946_ (.I(_04194_),
    .Z(_00644_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08947_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[22][15] ),
    .I1(_04054_),
    .S(_04189_),
    .Z(_04195_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08948_ (.I(_04195_),
    .Z(_00645_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08949_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[22][16] ),
    .I1(_02335_),
    .S(_04189_),
    .Z(_04196_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08950_ (.I(_04196_),
    .Z(_00646_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08951_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[22][17] ),
    .I1(_02337_),
    .S(_04189_),
    .Z(_04197_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08952_ (.I(_04197_),
    .Z(_00647_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08953_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[22][18] ),
    .I1(_02339_),
    .S(_04189_),
    .Z(_04198_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08954_ (.I(_04198_),
    .Z(_00648_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08955_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[22][19] ),
    .I1(_02341_),
    .S(_04189_),
    .Z(_04199_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08956_ (.I(_04199_),
    .Z(_00649_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08957_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[22][20] ),
    .I1(_02343_),
    .S(_04177_),
    .Z(_04200_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08958_ (.I(_04200_),
    .Z(_00650_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08959_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[22][21] ),
    .I1(_04061_),
    .S(_04177_),
    .Z(_04201_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08960_ (.I(_04201_),
    .Z(_00651_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08961_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[22][22] ),
    .I1(_04063_),
    .S(_04177_),
    .Z(_04202_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08962_ (.I(_04202_),
    .Z(_00652_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08963_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[22][23] ),
    .I1(_04065_),
    .S(_04177_),
    .Z(_04203_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08964_ (.I(_04203_),
    .Z(_00653_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08965_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[22][24] ),
    .I1(_04067_),
    .S(_04177_),
    .Z(_04204_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08966_ (.I(_04204_),
    .Z(_00654_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08967_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[22][25] ),
    .I1(_04069_),
    .S(_04177_),
    .Z(_04205_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08968_ (.I(_04205_),
    .Z(_00655_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08969_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[22][26] ),
    .I1(_03927_),
    .S(_04177_),
    .Z(_04206_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08970_ (.I(_04206_),
    .Z(_00656_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08971_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[22][27] ),
    .I1(_02351_),
    .S(_04177_),
    .Z(_04207_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08972_ (.I(_04207_),
    .Z(_00657_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08973_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[22][28] ),
    .I1(_02353_),
    .S(_04177_),
    .Z(_04208_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08974_ (.I(_04208_),
    .Z(_00658_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _08975_ (.A1(_02311_),
    .A2(_04175_),
    .ZN(_04209_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _08976_ (.I(_04209_),
    .Z(_04210_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08977_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[21][0] ),
    .I1(_02310_),
    .S(_04210_),
    .Z(_04211_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08978_ (.I(_04211_),
    .Z(_00659_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08979_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[21][1] ),
    .I1(_02393_),
    .S(_04210_),
    .Z(_04212_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08980_ (.I(_04212_),
    .Z(_00660_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08981_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[21][2] ),
    .I1(_02395_),
    .S(_04210_),
    .Z(_04213_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08982_ (.I(_04213_),
    .Z(_00661_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08983_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[21][3] ),
    .I1(_02397_),
    .S(_04210_),
    .Z(_04214_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08984_ (.I(_04214_),
    .Z(_00662_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08985_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[21][4] ),
    .I1(_02399_),
    .S(_04210_),
    .Z(_04215_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08986_ (.I(_04215_),
    .Z(_00663_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08987_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[21][5] ),
    .I1(_02401_),
    .S(_04210_),
    .Z(_04216_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08988_ (.I(_04216_),
    .Z(_00664_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08989_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[21][6] ),
    .I1(_02403_),
    .S(_04210_),
    .Z(_04217_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08990_ (.I(_04217_),
    .Z(_00665_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08991_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[21][7] ),
    .I1(_02405_),
    .S(_04210_),
    .Z(_04218_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08992_ (.I(_04218_),
    .Z(_00666_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08993_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[21][8] ),
    .I1(_02407_),
    .S(_04210_),
    .Z(_04219_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08994_ (.I(_04219_),
    .Z(_00667_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08995_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[21][9] ),
    .I1(_02409_),
    .S(_04210_),
    .Z(_04220_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08996_ (.I(_04220_),
    .Z(_00668_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _08997_ (.I(_04209_),
    .Z(_04221_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08998_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[21][10] ),
    .I1(_02411_),
    .S(_04221_),
    .Z(_04222_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08999_ (.I(_04222_),
    .Z(_00669_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09000_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[21][11] ),
    .I1(_02414_),
    .S(_04221_),
    .Z(_04223_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09001_ (.I(_04223_),
    .Z(_00670_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09002_ (.I(_04221_),
    .Z(_04224_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09003_ (.I(_04209_),
    .Z(_04225_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09004_ (.A1(_04047_),
    .A2(_04225_),
    .ZN(_04226_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09005_ (.A1(_03112_),
    .A2(_04224_),
    .B(_04226_),
    .ZN(_00671_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09006_ (.A1(_04050_),
    .A2(_04225_),
    .ZN(_04227_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09007_ (.A1(_03189_),
    .A2(_04224_),
    .B(_04227_),
    .ZN(_00672_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09008_ (.A1(_04052_),
    .A2(_04225_),
    .ZN(_04228_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09009_ (.A1(_03291_),
    .A2(_04224_),
    .B(_04228_),
    .ZN(_00673_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09010_ (.A1(_04054_),
    .A2(_04225_),
    .ZN(_04229_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09011_ (.A1(_03387_),
    .A2(_04224_),
    .B(_04229_),
    .ZN(_00674_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09012_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[21][16] ),
    .I1(_02335_),
    .S(_04221_),
    .Z(_04230_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09013_ (.I(_04230_),
    .Z(_00675_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09014_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[21][17] ),
    .I1(_02337_),
    .S(_04221_),
    .Z(_04231_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09015_ (.I(_04231_),
    .Z(_00676_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09016_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[21][18] ),
    .I1(_02339_),
    .S(_04221_),
    .Z(_04232_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09017_ (.I(_04232_),
    .Z(_00677_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09018_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[21][19] ),
    .I1(_02341_),
    .S(_04221_),
    .Z(_04233_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09019_ (.I(_04233_),
    .Z(_00678_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09020_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[21][20] ),
    .I1(_02343_),
    .S(_04221_),
    .Z(_04234_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09021_ (.I(_04234_),
    .Z(_00679_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09022_ (.A1(_04061_),
    .A2(_04225_),
    .ZN(_04235_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09023_ (.A1(_03557_),
    .A2(_04224_),
    .B(_04235_),
    .ZN(_00680_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09024_ (.A1(_04063_),
    .A2(_04225_),
    .ZN(_04236_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09025_ (.A1(_03485_),
    .A2(_04224_),
    .B(_04236_),
    .ZN(_00681_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09026_ (.A1(_04065_),
    .A2(_04225_),
    .ZN(_04237_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09027_ (.A1(_03434_),
    .A2(_04224_),
    .B(_04237_),
    .ZN(_00682_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09028_ (.A1(_04067_),
    .A2(_04225_),
    .ZN(_04238_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09029_ (.A1(_03338_),
    .A2(_04224_),
    .B(_04238_),
    .ZN(_00683_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09030_ (.A1(_04069_),
    .A2(_04225_),
    .ZN(_04239_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09031_ (.A1(_03240_),
    .A2(_04224_),
    .B(_04239_),
    .ZN(_00684_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09032_ (.A1(_03927_),
    .A2(_04225_),
    .ZN(_04240_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09033_ (.A1(_03148_),
    .A2(_04224_),
    .B(_04240_),
    .ZN(_00685_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09034_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[21][27] ),
    .I1(_02351_),
    .S(_04221_),
    .Z(_04241_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09035_ (.I(_04241_),
    .Z(_00686_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09036_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[21][28] ),
    .I1(_02353_),
    .S(_04221_),
    .Z(_04242_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09037_ (.I(_04242_),
    .Z(_00687_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09038_ (.I(_01378_),
    .Z(_04243_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09039_ (.I(_01408_),
    .ZN(_04244_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09040_ (.A1(\soc.spi_video_ram_1.fifo_read_request ),
    .A2(_04244_),
    .B(\soc.spi_video_ram_1.write_fifo.read_pointer[0] ),
    .ZN(_04245_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _09041_ (.A1(\soc.spi_video_ram_1.write_fifo.read_pointer[0] ),
    .A2(\soc.spi_video_ram_1.fifo_read_request ),
    .A3(_04244_),
    .Z(_04246_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _09042_ (.A1(_04243_),
    .A2(_04245_),
    .A3(_04246_),
    .ZN(_00688_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09043_ (.A1(\soc.spi_video_ram_1.write_fifo.read_pointer[1] ),
    .A2(_04246_),
    .Z(_04247_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09044_ (.I(_01379_),
    .Z(_04248_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09045_ (.A1(\soc.spi_video_ram_1.write_fifo.read_pointer[1] ),
    .A2(_04246_),
    .B(_04248_),
    .ZN(_04249_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09046_ (.A1(_04247_),
    .A2(_04249_),
    .ZN(_00689_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09047_ (.A1(\soc.spi_video_ram_1.write_fifo.read_pointer[2] ),
    .A2(_04247_),
    .ZN(_04250_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09048_ (.A1(\soc.spi_video_ram_1.write_fifo.read_pointer[2] ),
    .A2(_04247_),
    .Z(_04251_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _09049_ (.A1(_04243_),
    .A2(_04250_),
    .A3(_04251_),
    .ZN(_00690_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09050_ (.A1(\soc.spi_video_ram_1.write_fifo.read_pointer[3] ),
    .A2(_04251_),
    .ZN(_04252_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09051_ (.A1(\soc.spi_video_ram_1.write_fifo.read_pointer[3] ),
    .A2(_04251_),
    .Z(_04253_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _09052_ (.A1(_04243_),
    .A2(_04252_),
    .A3(_04253_),
    .ZN(_00691_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09053_ (.I(_01380_),
    .Z(_04254_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09054_ (.A1(\soc.spi_video_ram_1.write_fifo.read_pointer[4] ),
    .A2(_04253_),
    .Z(_04255_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09055_ (.A1(_04254_),
    .A2(_04255_),
    .Z(_04256_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09056_ (.I(_04256_),
    .Z(_00692_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _09057_ (.A1(_02116_),
    .A2(_04107_),
    .A3(_02214_),
    .ZN(_04257_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _09058_ (.I(_04257_),
    .Z(_04258_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _09059_ (.I(_04258_),
    .Z(_04259_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09060_ (.I0(_02213_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[20][0] ),
    .S(_04259_),
    .Z(_04260_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09061_ (.I(_04260_),
    .Z(_00693_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09062_ (.I0(_02219_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[20][1] ),
    .S(_04259_),
    .Z(_04261_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09063_ (.I(_04261_),
    .Z(_00694_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09064_ (.I0(_02221_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[20][2] ),
    .S(_04259_),
    .Z(_04262_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09065_ (.I(_04262_),
    .Z(_00695_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09066_ (.I0(_02223_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[20][3] ),
    .S(_04259_),
    .Z(_04263_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09067_ (.I(_04263_),
    .Z(_00696_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09068_ (.I0(_02225_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[20][4] ),
    .S(_04259_),
    .Z(_04264_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09069_ (.I(_04264_),
    .Z(_00697_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09070_ (.I0(_02227_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[20][5] ),
    .S(_04259_),
    .Z(_04265_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09071_ (.I(_04265_),
    .Z(_00698_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09072_ (.I0(_02229_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[20][6] ),
    .S(_04259_),
    .Z(_04266_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09073_ (.I(_04266_),
    .Z(_00699_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09074_ (.I0(_02231_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[20][7] ),
    .S(_04259_),
    .Z(_04267_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09075_ (.I(_04267_),
    .Z(_00700_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09076_ (.I0(_02233_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[20][8] ),
    .S(_04259_),
    .Z(_04268_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09077_ (.I(_04268_),
    .Z(_00701_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09078_ (.I0(_02235_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[20][9] ),
    .S(_04259_),
    .Z(_04269_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09079_ (.I(_04269_),
    .Z(_00702_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _09080_ (.I(_04257_),
    .Z(_04270_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09081_ (.I0(_02237_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[20][10] ),
    .S(_04270_),
    .Z(_04271_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09082_ (.I(_04271_),
    .Z(_00703_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09083_ (.I0(_02240_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[20][11] ),
    .S(_04270_),
    .Z(_04272_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09084_ (.I(_04272_),
    .Z(_00704_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09085_ (.I0(_02145_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[20][12] ),
    .S(_04270_),
    .Z(_04273_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09086_ (.I(_04273_),
    .Z(_00705_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09087_ (.I0(_02244_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[20][13] ),
    .S(_04270_),
    .Z(_04274_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09088_ (.I(_04274_),
    .Z(_00706_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09089_ (.I0(_02246_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[20][14] ),
    .S(_04270_),
    .Z(_04275_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09090_ (.I(_04275_),
    .Z(_00707_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09091_ (.I0(_02248_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[20][15] ),
    .S(_04270_),
    .Z(_04276_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09092_ (.I(_04276_),
    .Z(_00708_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09093_ (.I0(_02250_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[20][16] ),
    .S(_04270_),
    .Z(_04277_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09094_ (.I(_04277_),
    .Z(_00709_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09095_ (.I0(_02252_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[20][17] ),
    .S(_04270_),
    .Z(_04278_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09096_ (.I(_04278_),
    .Z(_00710_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09097_ (.I0(_02254_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[20][18] ),
    .S(_04270_),
    .Z(_04279_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09098_ (.I(_04279_),
    .Z(_00711_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09099_ (.I0(_02256_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[20][19] ),
    .S(_04270_),
    .Z(_04280_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09100_ (.I(_04280_),
    .Z(_00712_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09101_ (.I0(_02258_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[20][20] ),
    .S(_04258_),
    .Z(_04281_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09102_ (.I(_04281_),
    .Z(_00713_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09103_ (.I0(_02163_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[20][21] ),
    .S(_04258_),
    .Z(_04282_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09104_ (.I(_04282_),
    .Z(_00714_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09105_ (.I0(_02165_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[20][22] ),
    .S(_04258_),
    .Z(_04283_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09106_ (.I(_04283_),
    .Z(_00715_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09107_ (.I0(_02167_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[20][23] ),
    .S(_04258_),
    .Z(_04284_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09108_ (.I(_04284_),
    .Z(_00716_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09109_ (.I0(_02169_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[20][24] ),
    .S(_04258_),
    .Z(_04285_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09110_ (.I(_04285_),
    .Z(_00717_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09111_ (.I0(_02171_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[20][25] ),
    .S(_04258_),
    .Z(_04286_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09112_ (.I(_04286_),
    .Z(_00718_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09113_ (.I0(_02173_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[20][26] ),
    .S(_04258_),
    .Z(_04287_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09114_ (.I(_04287_),
    .Z(_00719_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09115_ (.I0(_02272_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[20][27] ),
    .S(_04258_),
    .Z(_04288_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09116_ (.I(_04288_),
    .Z(_00720_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09117_ (.I0(_02274_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[20][28] ),
    .S(_04258_),
    .Z(_04289_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09118_ (.I(_04289_),
    .Z(_00721_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09119_ (.I(\soc.spi_video_ram_1.current_state[2] ),
    .ZN(_04290_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09120_ (.A1(_04290_),
    .A2(_02673_),
    .B1(_01434_),
    .B2(_01419_),
    .ZN(_04291_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _09121_ (.A1(_01394_),
    .A2(_01429_),
    .A3(_01438_),
    .A4(_04291_),
    .ZN(_04292_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09122_ (.A1(_01414_),
    .A2(_04292_),
    .B(_01379_),
    .ZN(_04293_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09123_ (.I(_04293_),
    .Z(_04294_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09124_ (.A1(\soc.spi_video_ram_1.state_counter[0] ),
    .A2(_04294_),
    .ZN(_00722_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09125_ (.A1(\soc.spi_video_ram_1.state_counter[1] ),
    .A2(\soc.spi_video_ram_1.state_counter[0] ),
    .ZN(_04295_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09126_ (.A1(_04294_),
    .A2(_04295_),
    .ZN(_00723_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _09127_ (.A1(\soc.spi_video_ram_1.state_counter[1] ),
    .A2(\soc.spi_video_ram_1.state_counter[0] ),
    .A3(\soc.spi_video_ram_1.state_counter[2] ),
    .Z(_04296_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09128_ (.A1(\soc.spi_video_ram_1.state_counter[1] ),
    .A2(\soc.spi_video_ram_1.state_counter[0] ),
    .B(\soc.spi_video_ram_1.state_counter[2] ),
    .ZN(_04297_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _09129_ (.A1(_04294_),
    .A2(_04296_),
    .A3(_04297_),
    .ZN(_00724_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09130_ (.A1(\soc.spi_video_ram_1.state_counter[3] ),
    .A2(_04296_),
    .Z(_04298_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09131_ (.A1(\soc.spi_video_ram_1.state_counter[3] ),
    .A2(_04296_),
    .ZN(_04299_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _09132_ (.A1(_04294_),
    .A2(_04298_),
    .A3(_04299_),
    .ZN(_00725_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09133_ (.A1(\soc.spi_video_ram_1.state_counter[4] ),
    .A2(_04298_),
    .Z(_04300_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09134_ (.A1(\soc.spi_video_ram_1.state_counter[4] ),
    .A2(_04298_),
    .ZN(_04301_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _09135_ (.A1(_04294_),
    .A2(_04300_),
    .A3(_04301_),
    .ZN(_00726_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09136_ (.A1(\soc.spi_video_ram_1.state_counter[5] ),
    .A2(_04300_),
    .Z(_04302_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09137_ (.A1(\soc.spi_video_ram_1.state_counter[5] ),
    .A2(_04300_),
    .ZN(_04303_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _09138_ (.A1(_04294_),
    .A2(_04302_),
    .A3(_04303_),
    .ZN(_00727_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09139_ (.A1(\soc.spi_video_ram_1.state_counter[6] ),
    .A2(_04302_),
    .Z(_04304_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09140_ (.A1(\soc.spi_video_ram_1.state_counter[6] ),
    .A2(_04302_),
    .ZN(_04305_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _09141_ (.A1(_04294_),
    .A2(_04304_),
    .A3(_04305_),
    .ZN(_00728_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09142_ (.A1(\soc.spi_video_ram_1.state_counter[7] ),
    .A2(_04304_),
    .Z(_04306_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09143_ (.A1(\soc.spi_video_ram_1.state_counter[7] ),
    .A2(_04304_),
    .ZN(_04307_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _09144_ (.A1(_04294_),
    .A2(_04306_),
    .A3(_04307_),
    .ZN(_00729_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09145_ (.A1(\soc.spi_video_ram_1.state_counter[8] ),
    .A2(_04306_),
    .Z(_04308_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09146_ (.A1(\soc.spi_video_ram_1.state_counter[8] ),
    .A2(_04306_),
    .ZN(_04309_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _09147_ (.A1(_04293_),
    .A2(_04308_),
    .A3(_04309_),
    .ZN(_00730_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09148_ (.A1(\soc.spi_video_ram_1.state_counter[9] ),
    .A2(_04308_),
    .ZN(_04310_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09149_ (.A1(_04294_),
    .A2(_04310_),
    .ZN(_00731_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09150_ (.A1(\soc.spi_video_ram_1.state_counter[9] ),
    .A2(_04308_),
    .ZN(_04311_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09151_ (.A1(\soc.spi_video_ram_1.state_counter[10] ),
    .A2(_04311_),
    .Z(_04312_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09152_ (.A1(_04294_),
    .A2(_04312_),
    .ZN(_00732_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _09153_ (.A1(_01866_),
    .A2(_01959_),
    .A3(_03712_),
    .ZN(_04313_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _09154_ (.A1(_01860_),
    .A2(\soc.video_generator_1.v_count[8] ),
    .A3(\soc.video_generator_1.v_count[7] ),
    .A4(_01849_),
    .ZN(_04314_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _09155_ (.A1(_01931_),
    .A2(\soc.video_generator_1.v_count[1] ),
    .A3(_01866_),
    .ZN(_04315_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _09156_ (.A1(\soc.video_generator_1.v_count[2] ),
    .A2(_04314_),
    .A3(_04315_),
    .ZN(_04316_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_4 _09157_ (.A1(_01939_),
    .A2(_02034_),
    .A3(_04316_),
    .B(_01380_),
    .ZN(_04317_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09158_ (.A1(_01959_),
    .A2(_03712_),
    .ZN(_04318_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09159_ (.A1(\soc.video_generator_1.v_count[0] ),
    .A2(_04318_),
    .ZN(_04319_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _09160_ (.A1(_04313_),
    .A2(_04317_),
    .A3(_04319_),
    .ZN(_00733_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09161_ (.A1(\soc.video_generator_1.v_count[1] ),
    .A2(_04313_),
    .ZN(_04320_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09162_ (.A1(\soc.video_generator_1.v_count[1] ),
    .A2(_04313_),
    .Z(_04321_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _09163_ (.A1(_04317_),
    .A2(_04320_),
    .A3(_04321_),
    .ZN(_00734_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09164_ (.A1(\soc.video_generator_1.v_count[2] ),
    .A2(_04321_),
    .ZN(_04322_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09165_ (.A1(\soc.video_generator_1.v_count[2] ),
    .A2(_04321_),
    .Z(_04323_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _09166_ (.A1(_04317_),
    .A2(_04322_),
    .A3(_04323_),
    .ZN(_00735_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09167_ (.A1(\soc.video_generator_1.v_count[3] ),
    .A2(_04323_),
    .ZN(_04324_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09168_ (.A1(\soc.video_generator_1.v_count[3] ),
    .A2(_04323_),
    .Z(_04325_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _09169_ (.A1(_04317_),
    .A2(_04324_),
    .A3(_04325_),
    .ZN(_00736_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09170_ (.A1(_02034_),
    .A2(_04325_),
    .Z(_04326_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09171_ (.A1(_02034_),
    .A2(_04325_),
    .ZN(_04327_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _09172_ (.A1(_04317_),
    .A2(_04326_),
    .A3(_04327_),
    .ZN(_00737_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09173_ (.A1(_01939_),
    .A2(_02034_),
    .A3(_04325_),
    .ZN(_04328_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09174_ (.A1(_01939_),
    .A2(_04326_),
    .B(_04328_),
    .ZN(_04329_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09175_ (.A1(_04317_),
    .A2(_04329_),
    .ZN(_00738_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09176_ (.A1(_01849_),
    .A2(_04328_),
    .Z(_04330_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09177_ (.A1(_04317_),
    .A2(_04330_),
    .ZN(_00739_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09178_ (.I(\soc.video_generator_1.v_count[7] ),
    .ZN(_04331_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _09179_ (.A1(_01849_),
    .A2(_01939_),
    .A3(_02034_),
    .A4(_04325_),
    .ZN(_04332_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09180_ (.A1(_02034_),
    .A2(_04325_),
    .ZN(_04333_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09181_ (.A1(_01856_),
    .A2(_04333_),
    .ZN(_04334_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _09182_ (.A1(_04331_),
    .A2(_04332_),
    .B(_04334_),
    .C(_04317_),
    .ZN(_00740_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09183_ (.A1(\soc.video_generator_1.v_count[8] ),
    .A2(_04334_),
    .ZN(_04335_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09184_ (.A1(_01863_),
    .A2(_04333_),
    .ZN(_04336_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _09185_ (.A1(_04317_),
    .A2(_04335_),
    .A3(_04336_),
    .ZN(_00741_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09186_ (.A1(_01853_),
    .A2(_04336_),
    .ZN(_04337_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _09187_ (.A1(_01853_),
    .A2(_04336_),
    .B(_04337_),
    .C(_04317_),
    .ZN(_00742_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09188_ (.I(_01589_),
    .ZN(_04338_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _09189_ (.I(_01459_),
    .Z(_04339_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09190_ (.I0(_02213_),
    .I1(_04338_),
    .S(_04339_),
    .Z(_04340_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09191_ (.I(_04340_),
    .Z(_00743_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09192_ (.I(_01459_),
    .Z(_04341_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09193_ (.A1(\soc.spi_video_ram_1.fifo_in_data[1] ),
    .A2(_04341_),
    .ZN(_04342_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09194_ (.A1(_00011_),
    .A2(_01613_),
    .B(_04342_),
    .ZN(_00744_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09195_ (.A1(\soc.spi_video_ram_1.fifo_in_data[2] ),
    .A2(_04341_),
    .ZN(_04343_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09196_ (.A1(_00011_),
    .A2(_01632_),
    .B(_04343_),
    .ZN(_00745_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09197_ (.A1(\soc.spi_video_ram_1.fifo_in_data[3] ),
    .A2(_04341_),
    .ZN(_04344_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09198_ (.A1(_00011_),
    .A2(_01652_),
    .B(_04344_),
    .ZN(_00746_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09199_ (.A1(\soc.spi_video_ram_1.fifo_in_data[4] ),
    .A2(_04341_),
    .ZN(_04345_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09200_ (.A1(_00011_),
    .A2(_01666_),
    .B(_04345_),
    .ZN(_00747_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09201_ (.I(_01459_),
    .Z(_04346_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09202_ (.A1(\soc.spi_video_ram_1.fifo_in_data[5] ),
    .A2(_04346_),
    .ZN(_04347_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09203_ (.A1(_00011_),
    .A2(_01680_),
    .B(_04347_),
    .ZN(_00748_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09204_ (.A1(\soc.spi_video_ram_1.fifo_in_data[6] ),
    .A2(_04346_),
    .ZN(_04348_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09205_ (.A1(_00011_),
    .A2(_01699_),
    .B(_04348_),
    .ZN(_00749_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09206_ (.A1(\soc.spi_video_ram_1.fifo_in_data[7] ),
    .A2(_04346_),
    .ZN(_04349_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09207_ (.A1(_00011_),
    .A2(_01713_),
    .B(_04349_),
    .ZN(_00750_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09208_ (.A1(\soc.spi_video_ram_1.fifo_in_data[8] ),
    .A2(_04346_),
    .ZN(_04350_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09209_ (.A1(_00011_),
    .A2(_01736_),
    .B(_04350_),
    .ZN(_00751_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09210_ (.A1(\soc.spi_video_ram_1.fifo_in_data[9] ),
    .A2(_04346_),
    .ZN(_04351_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09211_ (.A1(_00011_),
    .A2(_01752_),
    .B(_04351_),
    .ZN(_00752_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09212_ (.A1(\soc.spi_video_ram_1.fifo_in_data[10] ),
    .A2(_04346_),
    .ZN(_04352_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09213_ (.A1(_04341_),
    .A2(_01767_),
    .B(_04352_),
    .ZN(_00753_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09214_ (.A1(\soc.spi_video_ram_1.fifo_in_data[11] ),
    .A2(_04346_),
    .ZN(_04353_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09215_ (.A1(_04341_),
    .A2(_01779_),
    .B(_04353_),
    .ZN(_00754_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09216_ (.A1(_04047_),
    .A2(_04346_),
    .ZN(_04354_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09217_ (.A1(_04341_),
    .A2(_01803_),
    .B(_04354_),
    .ZN(_00755_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09218_ (.A1(_04050_),
    .A2(_04346_),
    .ZN(_04355_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09219_ (.A1(_04341_),
    .A2(_01819_),
    .B(_04355_),
    .ZN(_00756_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09220_ (.A1(_04052_),
    .A2(_04346_),
    .ZN(_04356_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09221_ (.A1(_04341_),
    .A2(_01834_),
    .B(_04356_),
    .ZN(_00757_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09222_ (.A1(_04054_),
    .A2(_04339_),
    .ZN(_04357_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09223_ (.A1(_04341_),
    .A2(_02539_),
    .B(_04357_),
    .ZN(_00758_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09224_ (.A1(_02179_),
    .A2(_03729_),
    .ZN(_04358_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _09225_ (.I(_04358_),
    .Z(_04359_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 _09226_ (.I(_04359_),
    .Z(_04360_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09227_ (.I0(_02213_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[9][0] ),
    .S(_04360_),
    .Z(_04361_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09228_ (.I(_04361_),
    .Z(_00759_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09229_ (.I0(_02219_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[9][1] ),
    .S(_04360_),
    .Z(_04362_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09230_ (.I(_04362_),
    .Z(_00760_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09231_ (.I0(_02221_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[9][2] ),
    .S(_04360_),
    .Z(_04363_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09232_ (.I(_04363_),
    .Z(_00761_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09233_ (.I0(_02223_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[9][3] ),
    .S(_04360_),
    .Z(_04364_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09234_ (.I(_04364_),
    .Z(_00762_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _09235_ (.I(_04359_),
    .Z(_04365_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09236_ (.I0(_02225_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[9][4] ),
    .S(_04365_),
    .Z(_04366_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09237_ (.I(_04366_),
    .Z(_00763_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09238_ (.I0(_02227_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[9][5] ),
    .S(_04365_),
    .Z(_04367_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09239_ (.I(_04367_),
    .Z(_00764_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09240_ (.I0(_02229_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[9][6] ),
    .S(_04365_),
    .Z(_04368_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09241_ (.I(_04368_),
    .Z(_00765_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09242_ (.I0(_02231_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[9][7] ),
    .S(_04365_),
    .Z(_04369_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09243_ (.I(_04369_),
    .Z(_00766_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09244_ (.I0(_02233_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[9][8] ),
    .S(_04365_),
    .Z(_04370_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09245_ (.I(_04370_),
    .Z(_00767_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09246_ (.I0(_02235_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[9][9] ),
    .S(_04365_),
    .Z(_04371_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09247_ (.I(_04371_),
    .Z(_00768_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09248_ (.I0(_02237_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[9][10] ),
    .S(_04365_),
    .Z(_04372_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09249_ (.I(_04372_),
    .Z(_00769_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09250_ (.I0(_02240_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[9][11] ),
    .S(_04365_),
    .Z(_04373_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09251_ (.I(_04373_),
    .Z(_00770_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09252_ (.I0(_02242_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[9][12] ),
    .S(_04365_),
    .Z(_04374_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09253_ (.I(_04374_),
    .Z(_00771_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09254_ (.I(_04359_),
    .Z(_04375_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09255_ (.A1(_04050_),
    .A2(_04375_),
    .ZN(_04376_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09256_ (.A1(_03210_),
    .A2(_04375_),
    .B(_04376_),
    .ZN(_00772_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09257_ (.A1(_04052_),
    .A2(_04375_),
    .ZN(_04377_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09258_ (.A1(_03308_),
    .A2(_04375_),
    .B(_04377_),
    .ZN(_00773_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09259_ (.A1(_04054_),
    .A2(_04360_),
    .ZN(_04378_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09260_ (.A1(_03410_),
    .A2(_04375_),
    .B(_04378_),
    .ZN(_00774_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09261_ (.I0(_02250_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[9][16] ),
    .S(_04365_),
    .Z(_04379_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09262_ (.I(_04379_),
    .Z(_00775_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09263_ (.I0(_02252_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[9][17] ),
    .S(_04359_),
    .Z(_04380_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09264_ (.I(_04380_),
    .Z(_00776_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09265_ (.I0(_02254_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[9][18] ),
    .S(_04359_),
    .Z(_04381_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09266_ (.I(_04381_),
    .Z(_00777_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09267_ (.I0(_02256_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[9][19] ),
    .S(_04359_),
    .Z(_04382_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09268_ (.I(_04382_),
    .Z(_00778_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09269_ (.I0(_02258_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[9][20] ),
    .S(_04359_),
    .Z(_04383_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09270_ (.I(_04383_),
    .Z(_00779_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09271_ (.A1(_04061_),
    .A2(_04360_),
    .ZN(_04384_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09272_ (.A1(_03537_),
    .A2(_04375_),
    .B(_04384_),
    .ZN(_00780_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09273_ (.A1(_04063_),
    .A2(_04360_),
    .ZN(_04385_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09274_ (.A1(_03517_),
    .A2(_04375_),
    .B(_04385_),
    .ZN(_00781_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09275_ (.A1(_04065_),
    .A2(_04360_),
    .ZN(_04386_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09276_ (.A1(_03460_),
    .A2(_04375_),
    .B(_04386_),
    .ZN(_00782_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09277_ (.A1(_04067_),
    .A2(_04360_),
    .ZN(_04387_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09278_ (.A1(_03364_),
    .A2(_04375_),
    .B(_04387_),
    .ZN(_00783_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09279_ (.A1(_04069_),
    .A2(_04360_),
    .ZN(_04388_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09280_ (.A1(_03266_),
    .A2(_04375_),
    .B(_04388_),
    .ZN(_00784_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09281_ (.I0(_02270_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[9][26] ),
    .S(_04359_),
    .Z(_04389_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09282_ (.I(_04389_),
    .Z(_00785_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09283_ (.I0(_02272_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[9][27] ),
    .S(_04359_),
    .Z(_04390_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09284_ (.I(_04390_),
    .Z(_00786_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09285_ (.I0(_02274_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[9][28] ),
    .S(_04359_),
    .Z(_04391_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09286_ (.I(_04391_),
    .Z(_00787_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _09287_ (.A1(\soc.spi_video_ram_1.write_fifo.write_pointer[4] ),
    .A2(_01403_),
    .A3(_03862_),
    .ZN(_04392_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09288_ (.A1(_02214_),
    .A2(_04392_),
    .ZN(_04393_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _09289_ (.I(_04393_),
    .Z(_04394_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _09290_ (.I(_04394_),
    .Z(_04395_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09291_ (.I0(_02213_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[4][0] ),
    .S(_04395_),
    .Z(_04396_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09292_ (.I(_04396_),
    .Z(_00788_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09293_ (.I0(_02219_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[4][1] ),
    .S(_04395_),
    .Z(_04397_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09294_ (.I(_04397_),
    .Z(_00789_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09295_ (.I0(_02221_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[4][2] ),
    .S(_04395_),
    .Z(_04398_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09296_ (.I(_04398_),
    .Z(_00790_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09297_ (.I0(_02223_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[4][3] ),
    .S(_04395_),
    .Z(_04399_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09298_ (.I(_04399_),
    .Z(_00791_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09299_ (.I0(_02225_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[4][4] ),
    .S(_04395_),
    .Z(_04400_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09300_ (.I(_04400_),
    .Z(_00792_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09301_ (.I0(_02227_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[4][5] ),
    .S(_04395_),
    .Z(_04401_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09302_ (.I(_04401_),
    .Z(_00793_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09303_ (.I0(_02229_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[4][6] ),
    .S(_04395_),
    .Z(_04402_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09304_ (.I(_04402_),
    .Z(_00794_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09305_ (.I0(_02231_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[4][7] ),
    .S(_04395_),
    .Z(_04403_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09306_ (.I(_04403_),
    .Z(_00795_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09307_ (.I0(_02233_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[4][8] ),
    .S(_04395_),
    .Z(_04404_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09308_ (.I(_04404_),
    .Z(_00796_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09309_ (.I0(_02235_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[4][9] ),
    .S(_04395_),
    .Z(_04405_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09310_ (.I(_04405_),
    .Z(_00797_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _09311_ (.I(_04393_),
    .Z(_04406_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09312_ (.I0(_02237_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[4][10] ),
    .S(_04406_),
    .Z(_04407_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09313_ (.I(_04407_),
    .Z(_00798_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09314_ (.I0(_02240_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[4][11] ),
    .S(_04406_),
    .Z(_04408_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09315_ (.I(_04408_),
    .Z(_00799_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09316_ (.I0(_02242_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[4][12] ),
    .S(_04406_),
    .Z(_04409_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09317_ (.I(_04409_),
    .Z(_00800_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09318_ (.I0(_02244_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[4][13] ),
    .S(_04406_),
    .Z(_04410_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09319_ (.I(_04410_),
    .Z(_00801_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09320_ (.I0(_02246_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[4][14] ),
    .S(_04406_),
    .Z(_04411_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09321_ (.I(_04411_),
    .Z(_00802_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09322_ (.I0(_02248_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[4][15] ),
    .S(_04406_),
    .Z(_04412_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09323_ (.I(_04412_),
    .Z(_00803_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09324_ (.I0(_02250_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[4][16] ),
    .S(_04406_),
    .Z(_04413_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09325_ (.I(_04413_),
    .Z(_00804_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09326_ (.I0(_02252_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[4][17] ),
    .S(_04406_),
    .Z(_04414_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09327_ (.I(_04414_),
    .Z(_00805_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09328_ (.I0(_02254_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[4][18] ),
    .S(_04406_),
    .Z(_04415_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09329_ (.I(_04415_),
    .Z(_00806_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09330_ (.I0(_02256_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[4][19] ),
    .S(_04406_),
    .Z(_04416_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09331_ (.I(_04416_),
    .Z(_00807_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09332_ (.I0(_02258_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[4][20] ),
    .S(_04394_),
    .Z(_04417_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09333_ (.I(_04417_),
    .Z(_00808_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09334_ (.I0(_02260_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[4][21] ),
    .S(_04394_),
    .Z(_04418_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09335_ (.I(_04418_),
    .Z(_00809_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09336_ (.I0(_02262_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[4][22] ),
    .S(_04394_),
    .Z(_04419_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09337_ (.I(_04419_),
    .Z(_00810_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09338_ (.I0(_02264_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[4][23] ),
    .S(_04394_),
    .Z(_04420_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09339_ (.I(_04420_),
    .Z(_00811_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09340_ (.I0(_02266_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[4][24] ),
    .S(_04394_),
    .Z(_04421_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09341_ (.I(_04421_),
    .Z(_00812_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09342_ (.I0(_02268_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[4][25] ),
    .S(_04394_),
    .Z(_04422_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09343_ (.I(_04422_),
    .Z(_00813_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09344_ (.I0(_02270_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[4][26] ),
    .S(_04394_),
    .Z(_04423_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09345_ (.I(_04423_),
    .Z(_00814_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09346_ (.I0(_02272_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[4][27] ),
    .S(_04394_),
    .Z(_04424_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09347_ (.I(_04424_),
    .Z(_00815_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09348_ (.I0(_02274_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[4][28] ),
    .S(_04394_),
    .Z(_04425_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09349_ (.I(_04425_),
    .Z(_00816_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _09350_ (.I(\soc.rom_encoder_0.write_enable ),
    .ZN(_04426_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09351_ (.A1(_04426_),
    .A2(_01378_),
    .ZN(_04427_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09352_ (.I(_04427_),
    .Z(_00817_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _09353_ (.A1(\soc.spi_video_ram_1.current_state[3] ),
    .A2(\soc.spi_video_ram_1.current_state[1] ),
    .A3(\soc.spi_video_ram_1.current_state[0] ),
    .A4(\soc.spi_video_ram_1.current_state[2] ),
    .ZN(_04428_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09354_ (.A1(_04428_),
    .A2(_04295_),
    .ZN(_04429_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09355_ (.A1(\soc.spi_video_ram_1.state_counter[0] ),
    .A2(_04428_),
    .B(_04429_),
    .ZN(_04430_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09356_ (.A1(net69),
    .A2(_04430_),
    .ZN(_04431_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09357_ (.A1(\soc.spi_video_ram_1.state_sram_clk_counter[0] ),
    .A2(_04431_),
    .Z(_04432_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _09358_ (.A1(\soc.spi_video_ram_1.current_state[2] ),
    .A2(net68),
    .ZN(_04433_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09359_ (.A1(\soc.spi_video_ram_1.state_sram_clk_counter[0] ),
    .A2(_04431_),
    .B(_04433_),
    .ZN(_04434_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09360_ (.A1(_04432_),
    .A2(_04434_),
    .ZN(_00818_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09361_ (.A1(\soc.spi_video_ram_1.state_sram_clk_counter[1] ),
    .A2(_04432_),
    .Z(_04435_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09362_ (.A1(\soc.spi_video_ram_1.state_sram_clk_counter[1] ),
    .A2(_04432_),
    .B(_04433_),
    .ZN(_04436_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09363_ (.A1(_04435_),
    .A2(_04436_),
    .ZN(_00819_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09364_ (.A1(\soc.spi_video_ram_1.state_sram_clk_counter[2] ),
    .A2(_04435_),
    .Z(_04437_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09365_ (.A1(\soc.spi_video_ram_1.state_sram_clk_counter[2] ),
    .A2(_04435_),
    .B(_04433_),
    .ZN(_04438_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09366_ (.A1(_04437_),
    .A2(_04438_),
    .ZN(_00820_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09367_ (.A1(\soc.spi_video_ram_1.state_sram_clk_counter[3] ),
    .A2(_04437_),
    .Z(_04439_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09368_ (.A1(\soc.spi_video_ram_1.state_sram_clk_counter[3] ),
    .A2(_04437_),
    .B(_04433_),
    .ZN(_04440_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09369_ (.A1(_04439_),
    .A2(_04440_),
    .ZN(_00821_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09370_ (.A1(\soc.spi_video_ram_1.state_sram_clk_counter[4] ),
    .A2(_04439_),
    .Z(_04441_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09371_ (.A1(\soc.spi_video_ram_1.state_sram_clk_counter[4] ),
    .A2(_04439_),
    .B(_04433_),
    .ZN(_04442_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09372_ (.A1(_04441_),
    .A2(_04442_),
    .ZN(_00822_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09373_ (.A1(\soc.spi_video_ram_1.state_sram_clk_counter[5] ),
    .A2(_04441_),
    .Z(_04443_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09374_ (.A1(\soc.spi_video_ram_1.state_sram_clk_counter[5] ),
    .A2(_04441_),
    .B(_04433_),
    .ZN(_04444_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09375_ (.A1(_04443_),
    .A2(_04444_),
    .ZN(_00823_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09376_ (.A1(\soc.spi_video_ram_1.state_sram_clk_counter[6] ),
    .A2(_04443_),
    .Z(_04445_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09377_ (.A1(\soc.spi_video_ram_1.state_sram_clk_counter[6] ),
    .A2(_04443_),
    .B(_04433_),
    .ZN(_04446_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09378_ (.A1(_04445_),
    .A2(_04446_),
    .ZN(_00824_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09379_ (.A1(\soc.spi_video_ram_1.state_sram_clk_counter[7] ),
    .A2(_04445_),
    .B(_04433_),
    .ZN(_04447_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09380_ (.A1(\soc.spi_video_ram_1.state_sram_clk_counter[7] ),
    .A2(_04445_),
    .B(_04447_),
    .ZN(_00825_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _09381_ (.A1(\soc.spi_video_ram_1.current_state[2] ),
    .A2(net68),
    .Z(_04448_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09382_ (.A1(\soc.spi_video_ram_1.state_sram_clk_counter[7] ),
    .A2(_04445_),
    .ZN(_04449_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09383_ (.A1(_01387_),
    .A2(_04449_),
    .Z(_04450_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09384_ (.A1(_04448_),
    .A2(_04450_),
    .ZN(_00826_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09385_ (.A1(_04430_),
    .A2(_04448_),
    .ZN(_00827_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _09386_ (.A1(net69),
    .A2(_04430_),
    .A3(_04448_),
    .ZN(_00828_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _09387_ (.A1(net69),
    .A2(_04430_),
    .A3(_04433_),
    .Z(_04451_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09388_ (.I(_04451_),
    .Z(_00829_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09389_ (.A1(\soc.spi_video_ram_1.state_sram_clk_counter[2] ),
    .A2(\soc.spi_video_ram_1.state_sram_clk_counter[1] ),
    .B(\soc.spi_video_ram_1.state_sram_clk_counter[3] ),
    .ZN(_04452_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09390_ (.A1(_01388_),
    .A2(_04452_),
    .ZN(_04453_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _09391_ (.A1(_01387_),
    .A2(_04453_),
    .B(\soc.spi_video_ram_1.sram_sck_fall_edge ),
    .C(_01419_),
    .ZN(_04454_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09392_ (.I0(net9),
    .I1(\soc.spi_video_ram_1.read_value[0] ),
    .S(_04454_),
    .Z(_04455_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09393_ (.I(_04455_),
    .Z(_00831_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09394_ (.A1(net10),
    .A2(_04454_),
    .ZN(_04456_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09395_ (.A1(_02061_),
    .A2(_04454_),
    .B(_04456_),
    .ZN(_00832_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09396_ (.I0(net11),
    .I1(\soc.spi_video_ram_1.read_value[2] ),
    .S(_04454_),
    .Z(_04457_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09397_ (.I(_04457_),
    .Z(_00833_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09398_ (.I0(net12),
    .I1(\soc.spi_video_ram_1.read_value[3] ),
    .S(_04454_),
    .Z(_04458_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09399_ (.I(_04458_),
    .Z(_00834_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _09400_ (.A1(_02437_),
    .A2(_02447_),
    .ZN(_04459_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _09401_ (.A1(_04459_),
    .A2(_02460_),
    .B(_03765_),
    .C(_02445_),
    .ZN(_04460_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09402_ (.A1(\soc.rom_encoder_0.output_buffer[1] ),
    .A2(_04460_),
    .ZN(_04461_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09403_ (.A1(\soc.rom_encoder_0.output_buffer[5] ),
    .A2(_02541_),
    .ZN(_04462_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09404_ (.A1(\soc.rom_encoder_0.request_address[4] ),
    .A2(_02543_),
    .ZN(_04463_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _09405_ (.A1(_02542_),
    .A2(_04461_),
    .B(_04462_),
    .C(_04463_),
    .ZN(_00835_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09406_ (.A1(\soc.rom_encoder_0.output_buffer[2] ),
    .A2(_04460_),
    .ZN(_04464_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09407_ (.A1(\soc.rom_encoder_0.output_buffer[6] ),
    .A2(_02541_),
    .ZN(_04465_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09408_ (.A1(\soc.rom_encoder_0.request_address[5] ),
    .A2(_02543_),
    .ZN(_04466_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _09409_ (.A1(_02542_),
    .A2(_04464_),
    .B(_04465_),
    .C(_04466_),
    .ZN(_00836_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09410_ (.A1(\soc.rom_encoder_0.request_address[6] ),
    .A2(_02520_),
    .B(\soc.rom_encoder_0.output_buffer[3] ),
    .ZN(_04467_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09411_ (.I(\soc.rom_encoder_0.request_address[6] ),
    .ZN(_04468_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _09412_ (.A1(_04468_),
    .A2(_02441_),
    .B(_02515_),
    .C(_02454_),
    .ZN(_04469_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _09413_ (.A1(_02443_),
    .A2(_02441_),
    .B1(_04459_),
    .B2(_02460_),
    .C(_02445_),
    .ZN(_04470_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09414_ (.A1(_04469_),
    .A2(_04470_),
    .ZN(_04471_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09415_ (.A1(\soc.rom_encoder_0.output_buffer[7] ),
    .A2(_02541_),
    .ZN(_04472_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _09416_ (.A1(_02542_),
    .A2(_04467_),
    .A3(_04471_),
    .B(_04472_),
    .ZN(_00837_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09417_ (.I(_02541_),
    .Z(_04473_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09418_ (.A1(\soc.rom_encoder_0.request_data_out[0] ),
    .A2(_03767_),
    .Z(_04474_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _09419_ (.A1(\soc.rom_encoder_0.request_address[7] ),
    .A2(_02520_),
    .B1(_04460_),
    .B2(\soc.rom_encoder_0.output_buffer[4] ),
    .C(_04474_),
    .ZN(_04475_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09420_ (.A1(\soc.rom_encoder_0.output_buffer[8] ),
    .A2(_02542_),
    .ZN(_04476_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09421_ (.A1(_04473_),
    .A2(_04475_),
    .B(_04476_),
    .ZN(_00838_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09422_ (.A1(\soc.rom_encoder_0.request_data_out[1] ),
    .A2(_03767_),
    .Z(_04477_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _09423_ (.A1(\soc.rom_encoder_0.request_address[8] ),
    .A2(_02520_),
    .B1(_04460_),
    .B2(\soc.rom_encoder_0.output_buffer[5] ),
    .C(_04477_),
    .ZN(_04478_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09424_ (.I(_02541_),
    .Z(_04479_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09425_ (.A1(\soc.rom_encoder_0.output_buffer[9] ),
    .A2(_04479_),
    .ZN(_04480_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09426_ (.A1(_04473_),
    .A2(_04478_),
    .B(_04480_),
    .ZN(_00839_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09427_ (.A1(\soc.rom_encoder_0.request_data_out[2] ),
    .A2(_03767_),
    .Z(_04481_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _09428_ (.A1(\soc.rom_encoder_0.request_address[9] ),
    .A2(_02520_),
    .B1(_04460_),
    .B2(\soc.rom_encoder_0.output_buffer[6] ),
    .C(_04481_),
    .ZN(_04482_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09429_ (.A1(\soc.rom_encoder_0.output_buffer[10] ),
    .A2(_04479_),
    .ZN(_04483_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09430_ (.A1(_04473_),
    .A2(_04482_),
    .B(_04483_),
    .ZN(_00840_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09431_ (.A1(\soc.rom_encoder_0.request_data_out[3] ),
    .A2(_03767_),
    .Z(_04484_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _09432_ (.A1(\soc.rom_encoder_0.request_address[10] ),
    .A2(_02520_),
    .B1(_04460_),
    .B2(\soc.rom_encoder_0.output_buffer[7] ),
    .C(_04484_),
    .ZN(_04485_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09433_ (.A1(\soc.rom_encoder_0.output_buffer[11] ),
    .A2(_04479_),
    .ZN(_04486_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09434_ (.A1(_04473_),
    .A2(_04485_),
    .B(_04486_),
    .ZN(_00841_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09435_ (.A1(\soc.rom_encoder_0.request_data_out[4] ),
    .A2(_03767_),
    .Z(_04487_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _09436_ (.A1(\soc.rom_encoder_0.request_address[11] ),
    .A2(_02520_),
    .B1(_04460_),
    .B2(\soc.rom_encoder_0.output_buffer[8] ),
    .C(_04487_),
    .ZN(_04488_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09437_ (.A1(\soc.rom_encoder_0.output_buffer[12] ),
    .A2(_04479_),
    .ZN(_04489_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09438_ (.A1(_04473_),
    .A2(_04488_),
    .B(_04489_),
    .ZN(_00842_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09439_ (.A1(\soc.rom_encoder_0.request_data_out[5] ),
    .A2(_03767_),
    .Z(_04490_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _09440_ (.A1(\soc.rom_encoder_0.request_address[12] ),
    .A2(_02520_),
    .B1(_04460_),
    .B2(\soc.rom_encoder_0.output_buffer[9] ),
    .C(_04490_),
    .ZN(_04491_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09441_ (.A1(\soc.rom_encoder_0.output_buffer[13] ),
    .A2(_04479_),
    .ZN(_04492_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09442_ (.A1(_04473_),
    .A2(_04491_),
    .B(_04492_),
    .ZN(_00843_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09443_ (.A1(\soc.rom_encoder_0.request_data_out[6] ),
    .A2(_03767_),
    .Z(_04493_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _09444_ (.A1(\soc.rom_encoder_0.request_address[13] ),
    .A2(_02520_),
    .B1(_04460_),
    .B2(\soc.rom_encoder_0.output_buffer[10] ),
    .C(_04493_),
    .ZN(_04494_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09445_ (.A1(\soc.rom_encoder_0.output_buffer[14] ),
    .A2(_04479_),
    .ZN(_04495_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09446_ (.A1(_04473_),
    .A2(_04494_),
    .B(_04495_),
    .ZN(_00844_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09447_ (.A1(\soc.rom_encoder_0.request_data_out[7] ),
    .A2(_03767_),
    .Z(_04496_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _09448_ (.A1(\soc.rom_encoder_0.request_address[14] ),
    .A2(_02520_),
    .B1(_04460_),
    .B2(\soc.rom_encoder_0.output_buffer[11] ),
    .C(_04496_),
    .ZN(_04497_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09449_ (.A1(\soc.rom_encoder_0.output_buffer[15] ),
    .A2(_04479_),
    .ZN(_04498_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09450_ (.A1(_04473_),
    .A2(_04497_),
    .B(_04498_),
    .ZN(_00845_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09451_ (.I(\soc.rom_encoder_0.request_write ),
    .ZN(_04499_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09452_ (.A1(_04499_),
    .A2(_02525_),
    .B1(_03767_),
    .B2(\soc.rom_encoder_0.request_data_out[8] ),
    .ZN(_04500_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09453_ (.A1(_02458_),
    .A2(_03766_),
    .B(\soc.rom_encoder_0.output_buffer[12] ),
    .ZN(_04501_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09454_ (.A1(_04500_),
    .A2(_04501_),
    .ZN(_04502_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _09455_ (.A1(_02461_),
    .A2(_02541_),
    .A3(_04502_),
    .ZN(_04503_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09456_ (.A1(_03770_),
    .A2(_04473_),
    .B(_04503_),
    .ZN(_00846_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09457_ (.A1(_02445_),
    .A2(_02441_),
    .A3(_04459_),
    .ZN(_04504_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09458_ (.A1(\soc.rom_encoder_0.request_data_out[9] ),
    .A2(_02441_),
    .ZN(_04505_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09459_ (.A1(_02435_),
    .A2(_04505_),
    .B(_02524_),
    .ZN(_04506_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _09460_ (.A1(\soc.rom_encoder_0.output_buffer[13] ),
    .A2(_04504_),
    .B(_04506_),
    .C(_02461_),
    .ZN(_04507_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09461_ (.A1(\soc.rom_encoder_0.output_buffer[17] ),
    .A2(_04479_),
    .ZN(_04508_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09462_ (.A1(_04473_),
    .A2(_04507_),
    .B(_04508_),
    .ZN(_00847_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09463_ (.A1(\soc.rom_encoder_0.output_buffer[14] ),
    .A2(_02463_),
    .B1(_02464_),
    .B2(\soc.rom_encoder_0.request_data_out[10] ),
    .ZN(_04509_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09464_ (.A1(_02443_),
    .A2(_04509_),
    .ZN(_04510_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _09465_ (.A1(\soc.rom_encoder_0.output_buffer[14] ),
    .A2(_02455_),
    .B(_04510_),
    .C(_02461_),
    .ZN(_04511_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09466_ (.A1(\soc.rom_encoder_0.output_buffer[18] ),
    .A2(_04479_),
    .ZN(_04512_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09467_ (.A1(_02542_),
    .A2(_04511_),
    .B(_04512_),
    .ZN(_00848_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09468_ (.A1(\soc.rom_encoder_0.output_buffer[15] ),
    .A2(_02463_),
    .B1(_02464_),
    .B2(\soc.rom_encoder_0.request_data_out[11] ),
    .ZN(_04513_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09469_ (.A1(_02443_),
    .A2(_04513_),
    .ZN(_04514_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _09470_ (.A1(\soc.rom_encoder_0.output_buffer[15] ),
    .A2(_02455_),
    .B(_04514_),
    .C(_02461_),
    .ZN(_04515_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09471_ (.A1(\soc.rom_encoder_0.output_buffer[19] ),
    .A2(_04479_),
    .ZN(_04516_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09472_ (.A1(_02542_),
    .A2(_04515_),
    .B(_04516_),
    .ZN(_00849_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09473_ (.A1(_01437_),
    .A2(_01417_),
    .B(_02624_),
    .ZN(_04517_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09474_ (.A1(_01378_),
    .A2(_01410_),
    .ZN(_04518_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _09475_ (.A1(_02674_),
    .A2(_04517_),
    .B1(_04518_),
    .B2(_01392_),
    .ZN(_04519_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09476_ (.A1(_01379_),
    .A2(\soc.spi_video_ram_1.sram_sck_rise_edge ),
    .Z(_04520_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09477_ (.A1(_01428_),
    .A2(_04520_),
    .ZN(_04521_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09478_ (.A1(_01501_),
    .A2(_04521_),
    .Z(_04522_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09479_ (.A1(_04519_),
    .A2(_04522_),
    .ZN(_00850_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09480_ (.A1(_01501_),
    .A2(_04521_),
    .B(_01469_),
    .ZN(_04523_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _09481_ (.A1(_01485_),
    .A2(_04521_),
    .B(_04523_),
    .C(_04519_),
    .ZN(_00851_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09482_ (.A1(_01428_),
    .A2(_01485_),
    .ZN(_04524_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09483_ (.A1(_01518_),
    .A2(_04520_),
    .A3(_04524_),
    .ZN(_04525_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09484_ (.A1(_04520_),
    .A2(_04524_),
    .ZN(_04526_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09485_ (.A1(_01470_),
    .A2(_04526_),
    .ZN(_04527_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09486_ (.A1(_04519_),
    .A2(_04525_),
    .A3(_04527_),
    .ZN(_00852_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09487_ (.A1(_01463_),
    .A2(_04525_),
    .Z(_04528_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09488_ (.A1(_02882_),
    .A2(_04528_),
    .ZN(_00853_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09489_ (.A1(_01428_),
    .A2(_02091_),
    .ZN(_04529_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _09490_ (.A1(_01428_),
    .A2(_01465_),
    .B(_04520_),
    .C(_04529_),
    .ZN(_04530_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _09491_ (.A1(_01460_),
    .A2(_04520_),
    .B(_04530_),
    .C(_04519_),
    .ZN(_00854_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _09492_ (.A1(_01460_),
    .A2(_01464_),
    .A3(_04520_),
    .A4(_04524_),
    .ZN(_04531_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09493_ (.A1(\soc.spi_video_ram_1.buffer_index[5] ),
    .A2(_04531_),
    .Z(_04532_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09494_ (.A1(_02882_),
    .A2(_04532_),
    .ZN(_00855_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09495_ (.A1(_01387_),
    .A2(_04453_),
    .B(_01419_),
    .ZN(_00856_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09496_ (.I0(_02250_),
    .I1(\soc.cpu.AReg.data[0] ),
    .S(_04339_),
    .Z(_04533_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09497_ (.I(_04533_),
    .Z(_00857_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09498_ (.I0(_02252_),
    .I1(\soc.cpu.AReg.data[1] ),
    .S(_04339_),
    .Z(_04534_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09499_ (.I(_04534_),
    .Z(_00858_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09500_ (.I0(_02254_),
    .I1(\soc.cpu.AReg.data[2] ),
    .S(_04339_),
    .Z(_04535_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09501_ (.I(_04535_),
    .Z(_00859_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09502_ (.I0(_02256_),
    .I1(\soc.cpu.AReg.data[3] ),
    .S(_04339_),
    .Z(_04536_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09503_ (.I(_04536_),
    .Z(_00860_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09504_ (.I0(_02258_),
    .I1(\soc.cpu.AReg.data[4] ),
    .S(_04339_),
    .Z(_04537_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09505_ (.I(_04537_),
    .Z(_00861_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09506_ (.I0(_02260_),
    .I1(\soc.cpu.AReg.data[5] ),
    .S(_04339_),
    .Z(_04538_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09507_ (.I(_04538_),
    .Z(_00862_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09508_ (.I0(_02262_),
    .I1(\soc.cpu.AReg.data[6] ),
    .S(_04339_),
    .Z(_04539_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09509_ (.I(_04539_),
    .Z(_00863_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09510_ (.I0(_02264_),
    .I1(\soc.cpu.AReg.data[7] ),
    .S(_04339_),
    .Z(_04540_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09511_ (.I(_04540_),
    .Z(_00864_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09512_ (.I0(_02266_),
    .I1(\soc.cpu.AReg.data[8] ),
    .S(_01459_),
    .Z(_04541_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09513_ (.I(_04541_),
    .Z(_00865_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09514_ (.I0(_02268_),
    .I1(\soc.cpu.AReg.data[9] ),
    .S(_01459_),
    .Z(_04542_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09515_ (.I(_04542_),
    .Z(_00866_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09516_ (.I0(_02270_),
    .I1(\soc.cpu.AReg.data[10] ),
    .S(_01459_),
    .Z(_04543_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09517_ (.I(_04543_),
    .Z(_00867_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09518_ (.I0(_02272_),
    .I1(\soc.cpu.AReg.data[11] ),
    .S(_01459_),
    .Z(_04544_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09519_ (.I(_04544_),
    .Z(_00868_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09520_ (.I0(_02274_),
    .I1(\soc.cpu.AReg.data[12] ),
    .S(_01459_),
    .Z(_04545_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09521_ (.I(_04545_),
    .Z(_00869_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09522_ (.A1(_01994_),
    .A2(\soc.video_generator_1.h_count[4] ),
    .A3(\soc.video_generator_1.h_count[7] ),
    .ZN(_04546_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09523_ (.A1(\soc.spi_video_ram_1.initialized ),
    .A2(\soc.video_generator_1.h_count[1] ),
    .A3(_01839_),
    .ZN(_04547_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _09524_ (.A1(\soc.video_generator_1.h_count[6] ),
    .A2(_04546_),
    .A3(_04547_),
    .ZN(_04548_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _09525_ (.A1(_01836_),
    .A2(_01993_),
    .A3(_02058_),
    .A4(_04548_),
    .ZN(_04549_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09526_ (.A1(\soc.spi_video_ram_1.start_read ),
    .A2(_02673_),
    .ZN(_04550_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _09527_ (.A1(_02673_),
    .A2(_04549_),
    .B(_04550_),
    .C(_03714_),
    .ZN(_00870_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09528_ (.A1(_01430_),
    .A2(_01418_),
    .B(_01396_),
    .ZN(_00871_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09529_ (.I(_01451_),
    .ZN(_04551_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _09530_ (.A1(\soc.spi_video_ram_1.fifo_read_request ),
    .A2(_04551_),
    .B(\soc.spi_video_ram_1.fifo_write_request ),
    .ZN(_04552_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09531_ (.I(_01380_),
    .Z(_04553_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09532_ (.A1(_01444_),
    .A2(_04552_),
    .B(_04553_),
    .ZN(_04554_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09533_ (.A1(_01444_),
    .A2(_04552_),
    .B(_04554_),
    .ZN(_00872_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09534_ (.A1(_01441_),
    .A2(_04552_),
    .ZN(_04555_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09535_ (.A1(_01444_),
    .A2(_04552_),
    .ZN(_04556_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09536_ (.A1(\soc.spi_video_ram_1.write_fifo.write_pointer[1] ),
    .A2(_04556_),
    .B(_04254_),
    .ZN(_04557_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09537_ (.A1(_04555_),
    .A2(_04557_),
    .ZN(_00873_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09538_ (.A1(_01446_),
    .A2(_04552_),
    .ZN(_04558_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09539_ (.A1(_02116_),
    .A2(_04555_),
    .B(_04254_),
    .ZN(_04559_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09540_ (.A1(_04558_),
    .A2(_04559_),
    .ZN(_00874_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09541_ (.A1(_01446_),
    .A2(_04552_),
    .B(_02312_),
    .ZN(_04560_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09542_ (.A1(_01403_),
    .A2(_04558_),
    .ZN(_04561_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09543_ (.A1(_04254_),
    .A2(_04560_),
    .A3(_04561_),
    .ZN(_04562_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09544_ (.I(_04562_),
    .ZN(_00875_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09545_ (.A1(\soc.spi_video_ram_1.write_fifo.write_pointer[4] ),
    .A2(_04561_),
    .Z(_04563_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09546_ (.A1(_01396_),
    .A2(_04563_),
    .ZN(_00876_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _09547_ (.A1(_04243_),
    .A2(_04245_),
    .A3(_04246_),
    .ZN(_00877_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09548_ (.A1(_04247_),
    .A2(_04249_),
    .ZN(_00878_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _09549_ (.A1(_04243_),
    .A2(_04250_),
    .A3(_04251_),
    .ZN(_00879_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _09550_ (.A1(_04243_),
    .A2(_04252_),
    .A3(_04253_),
    .ZN(_00880_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09551_ (.A1(_04254_),
    .A2(_04255_),
    .Z(_04564_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09552_ (.I(_04564_),
    .Z(_00881_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09553_ (.A1(_02433_),
    .A2(_02442_),
    .Z(_04565_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _09554_ (.A1(_02434_),
    .A2(_02457_),
    .ZN(_04566_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09555_ (.A1(\soc.rom_encoder_0.current_state[2] ),
    .A2(_02447_),
    .ZN(_04567_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09556_ (.I(\soc.rom_encoder_0.input_bits_left[3] ),
    .ZN(_04568_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09557_ (.A1(\soc.rom_encoder_0.input_bits_left[2] ),
    .A2(_04568_),
    .ZN(_04569_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09558_ (.A1(\soc.rom_encoder_0.input_bits_left[4] ),
    .A2(_04569_),
    .ZN(_04570_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09559_ (.I(_04570_),
    .ZN(_04571_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09560_ (.A1(\soc.rom_encoder_0.request_write ),
    .A2(_02462_),
    .B(_04565_),
    .ZN(_04572_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _09561_ (.A1(_04567_),
    .A2(_04571_),
    .B(\soc.rom_encoder_0.toggled_sram_sck ),
    .C(_04572_),
    .ZN(_04573_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09562_ (.A1(_01378_),
    .A2(_04573_),
    .ZN(_04574_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09563_ (.A1(_04565_),
    .A2(_04566_),
    .B(_04574_),
    .ZN(_04575_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09564_ (.A1(\soc.rom_encoder_0.input_bits_left[2] ),
    .A2(_04575_),
    .ZN(_04576_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09565_ (.A1(\soc.rom_encoder_0.input_bits_left[2] ),
    .A2(_04575_),
    .ZN(_04577_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09566_ (.A1(\soc.rom_encoder_0.current_state[2] ),
    .A2(_04577_),
    .ZN(_04578_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09567_ (.A1(_04576_),
    .A2(_04578_),
    .ZN(_00882_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09568_ (.A1(_04565_),
    .A2(_04574_),
    .ZN(_04579_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09569_ (.A1(_04568_),
    .A2(_04577_),
    .ZN(_04580_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09570_ (.A1(\soc.rom_encoder_0.input_bits_left[2] ),
    .A2(_04575_),
    .B(\soc.rom_encoder_0.input_bits_left[3] ),
    .ZN(_04581_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09571_ (.A1(_04579_),
    .A2(_04580_),
    .A3(_04581_),
    .ZN(_00883_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09572_ (.A1(\soc.rom_encoder_0.input_bits_left[4] ),
    .A2(_04580_),
    .Z(_04582_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09573_ (.A1(_04579_),
    .A2(_04582_),
    .ZN(_00884_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09574_ (.I(\soc.rom_encoder_0.input_buffer[0] ),
    .ZN(_04583_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _09575_ (.A1(\soc.rom_encoder_0.toggled_sram_sck ),
    .A2(_04566_),
    .ZN(_04584_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09576_ (.I(_04584_),
    .Z(_04585_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09577_ (.I(_04584_),
    .Z(_04586_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09578_ (.A1(net5),
    .A2(_04586_),
    .B(_04553_),
    .ZN(_04587_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09579_ (.A1(_04583_),
    .A2(_04585_),
    .B(_04587_),
    .ZN(_00885_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09580_ (.I(\soc.rom_encoder_0.input_buffer[1] ),
    .ZN(_04588_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09581_ (.A1(net6),
    .A2(_04586_),
    .B(_04553_),
    .ZN(_04589_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09582_ (.A1(_04588_),
    .A2(_04585_),
    .B(_04589_),
    .ZN(_00886_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09583_ (.I(\soc.rom_encoder_0.input_buffer[2] ),
    .ZN(_04590_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09584_ (.A1(net7),
    .A2(_04586_),
    .B(_04553_),
    .ZN(_04591_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09585_ (.A1(_04590_),
    .A2(_04585_),
    .B(_04591_),
    .ZN(_00887_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09586_ (.I(\soc.rom_encoder_0.input_buffer[3] ),
    .ZN(_04592_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09587_ (.A1(net8),
    .A2(_04586_),
    .B(_04553_),
    .ZN(_04593_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09588_ (.A1(_04592_),
    .A2(_04585_),
    .B(_04593_),
    .ZN(_00888_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09589_ (.I(\soc.rom_encoder_0.input_buffer[4] ),
    .ZN(_04594_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09590_ (.A1(\soc.rom_encoder_0.input_buffer[0] ),
    .A2(_04586_),
    .B(_04553_),
    .ZN(_04595_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09591_ (.A1(_04594_),
    .A2(_04585_),
    .B(_04595_),
    .ZN(_00889_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09592_ (.I(\soc.rom_encoder_0.input_buffer[5] ),
    .ZN(_04596_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09593_ (.A1(\soc.rom_encoder_0.input_buffer[1] ),
    .A2(_04586_),
    .B(_04553_),
    .ZN(_04597_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09594_ (.A1(_04596_),
    .A2(_04585_),
    .B(_04597_),
    .ZN(_00890_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09595_ (.I(\soc.rom_encoder_0.input_buffer[6] ),
    .ZN(_04598_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09596_ (.A1(\soc.rom_encoder_0.input_buffer[2] ),
    .A2(_04586_),
    .B(_04553_),
    .ZN(_04599_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09597_ (.A1(_04598_),
    .A2(_04585_),
    .B(_04599_),
    .ZN(_00891_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09598_ (.I(\soc.rom_encoder_0.input_buffer[7] ),
    .ZN(_04600_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09599_ (.I(_01380_),
    .Z(_04601_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09600_ (.A1(\soc.rom_encoder_0.input_buffer[3] ),
    .A2(_04586_),
    .B(_04601_),
    .ZN(_04602_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09601_ (.A1(_04600_),
    .A2(_04585_),
    .B(_04602_),
    .ZN(_00892_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09602_ (.I(\soc.rom_encoder_0.input_buffer[8] ),
    .ZN(_04603_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09603_ (.A1(\soc.rom_encoder_0.input_buffer[4] ),
    .A2(_04584_),
    .B(_04601_),
    .ZN(_04604_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09604_ (.A1(_04603_),
    .A2(_04585_),
    .B(_04604_),
    .ZN(_00893_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09605_ (.I(\soc.rom_encoder_0.input_buffer[9] ),
    .ZN(_04605_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09606_ (.A1(\soc.rom_encoder_0.input_buffer[5] ),
    .A2(_04584_),
    .B(_04601_),
    .ZN(_04606_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09607_ (.A1(_04605_),
    .A2(_04585_),
    .B(_04606_),
    .ZN(_00894_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09608_ (.I(\soc.rom_encoder_0.input_buffer[10] ),
    .ZN(_04607_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09609_ (.A1(\soc.rom_encoder_0.input_buffer[6] ),
    .A2(_04584_),
    .B(_04601_),
    .ZN(_04608_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09610_ (.A1(_04607_),
    .A2(_04586_),
    .B(_04608_),
    .ZN(_00895_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09611_ (.I(\soc.rom_encoder_0.input_buffer[11] ),
    .ZN(_04609_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09612_ (.A1(\soc.rom_encoder_0.input_buffer[7] ),
    .A2(_04584_),
    .B(_04601_),
    .ZN(_04610_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09613_ (.A1(_04609_),
    .A2(_04586_),
    .B(_04610_),
    .ZN(_00896_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09614_ (.A1(\soc.rom_encoder_0.current_state[2] ),
    .A2(_02457_),
    .ZN(_04611_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09615_ (.A1(_02434_),
    .A2(_02447_),
    .ZN(_04612_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09616_ (.I0(\soc.hack_rom_request ),
    .I1(\soc.rom_loader.rom_request ),
    .S(\soc.rom_encoder_0.write_enable ),
    .Z(_04613_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09617_ (.A1(_04612_),
    .A2(_04613_),
    .B(\soc.rom_encoder_0.toggled_sram_sck ),
    .ZN(_04614_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _09618_ (.I(_04614_),
    .ZN(_04615_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09619_ (.A1(_01379_),
    .A2(_04611_),
    .A3(_04615_),
    .ZN(_04616_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _09620_ (.I(_04616_),
    .Z(_04617_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09621_ (.I(_04617_),
    .Z(_04618_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09622_ (.A1(\soc.rom_encoder_0.request_write ),
    .A2(_04618_),
    .ZN(_04619_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09623_ (.A1(_04426_),
    .A2(_04618_),
    .B(_04619_),
    .ZN(_00897_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09624_ (.I0(\soc.rom_encoder_0.data_out[0] ),
    .I1(\soc.rom_encoder_0.request_data_out[0] ),
    .S(_04618_),
    .Z(_04620_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09625_ (.I(_04620_),
    .Z(_00898_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _09626_ (.I(_04617_),
    .Z(_04621_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09627_ (.I0(\soc.rom_encoder_0.data_out[1] ),
    .I1(\soc.rom_encoder_0.request_data_out[1] ),
    .S(_04621_),
    .Z(_04622_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09628_ (.I(_04622_),
    .Z(_00899_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09629_ (.I0(\soc.rom_encoder_0.data_out[2] ),
    .I1(\soc.rom_encoder_0.request_data_out[2] ),
    .S(_04621_),
    .Z(_04623_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09630_ (.I(_04623_),
    .Z(_00900_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09631_ (.I0(\soc.rom_encoder_0.data_out[3] ),
    .I1(\soc.rom_encoder_0.request_data_out[3] ),
    .S(_04621_),
    .Z(_04624_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09632_ (.I(_04624_),
    .Z(_00901_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09633_ (.I0(\soc.rom_encoder_0.data_out[4] ),
    .I1(\soc.rom_encoder_0.request_data_out[4] ),
    .S(_04621_),
    .Z(_04625_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09634_ (.I(_04625_),
    .Z(_00902_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09635_ (.I0(\soc.rom_encoder_0.data_out[5] ),
    .I1(\soc.rom_encoder_0.request_data_out[5] ),
    .S(_04621_),
    .Z(_04626_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09636_ (.I(_04626_),
    .Z(_00903_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09637_ (.I0(\soc.rom_encoder_0.data_out[6] ),
    .I1(\soc.rom_encoder_0.request_data_out[6] ),
    .S(_04621_),
    .Z(_04627_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09638_ (.I(_04627_),
    .Z(_00904_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09639_ (.I0(\soc.rom_encoder_0.data_out[7] ),
    .I1(\soc.rom_encoder_0.request_data_out[7] ),
    .S(_04621_),
    .Z(_04628_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09640_ (.I(_04628_),
    .Z(_00905_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09641_ (.I0(\soc.rom_encoder_0.data_out[8] ),
    .I1(\soc.rom_encoder_0.request_data_out[8] ),
    .S(_04621_),
    .Z(_04629_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09642_ (.I(_04629_),
    .Z(_00906_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09643_ (.I0(\soc.rom_encoder_0.data_out[9] ),
    .I1(\soc.rom_encoder_0.request_data_out[9] ),
    .S(_04621_),
    .Z(_04630_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09644_ (.I(_04630_),
    .Z(_00907_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09645_ (.I0(\soc.rom_encoder_0.data_out[10] ),
    .I1(\soc.rom_encoder_0.request_data_out[10] ),
    .S(_04621_),
    .Z(_04631_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09646_ (.I(_04631_),
    .Z(_00908_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _09647_ (.I(_04617_),
    .Z(_04632_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09648_ (.I0(\soc.rom_encoder_0.data_out[11] ),
    .I1(\soc.rom_encoder_0.request_data_out[11] ),
    .S(_04632_),
    .Z(_04633_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09649_ (.I(_04633_),
    .Z(_00909_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09650_ (.I0(\soc.rom_encoder_0.data_out[12] ),
    .I1(\soc.rom_encoder_0.request_data_out[12] ),
    .S(_04632_),
    .Z(_04634_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09651_ (.I(_04634_),
    .Z(_00910_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09652_ (.I0(\soc.rom_encoder_0.data_out[13] ),
    .I1(\soc.rom_encoder_0.request_data_out[13] ),
    .S(_04632_),
    .Z(_04635_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09653_ (.I(_04635_),
    .Z(_00911_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09654_ (.I0(\soc.rom_encoder_0.data_out[14] ),
    .I1(\soc.rom_encoder_0.request_data_out[14] ),
    .S(_04632_),
    .Z(_04636_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09655_ (.I(_04636_),
    .Z(_00912_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09656_ (.I0(\soc.rom_encoder_0.data_out[15] ),
    .I1(\soc.rom_encoder_0.request_data_out[15] ),
    .S(_04632_),
    .Z(_04637_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09657_ (.I(_04637_),
    .Z(_00913_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _09658_ (.I(\soc.rom_encoder_0.write_enable ),
    .Z(_04638_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09659_ (.I(_04638_),
    .Z(_04639_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09660_ (.I0(\soc.cpu.PC.REG.data[0] ),
    .I1(\soc.rom_loader.current_address[0] ),
    .S(_04639_),
    .Z(_04640_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09661_ (.I0(_04640_),
    .I1(\soc.rom_encoder_0.request_address[0] ),
    .S(_04632_),
    .Z(_04641_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09662_ (.I(_04641_),
    .Z(_00914_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09663_ (.I0(\soc.cpu.PC.REG.data[1] ),
    .I1(\soc.rom_loader.current_address[1] ),
    .S(_04639_),
    .Z(_04642_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09664_ (.I0(_04642_),
    .I1(\soc.rom_encoder_0.request_address[1] ),
    .S(_04632_),
    .Z(_04643_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09665_ (.I(_04643_),
    .Z(_00915_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09666_ (.I0(\soc.cpu.PC.REG.data[2] ),
    .I1(\soc.rom_loader.current_address[2] ),
    .S(_04638_),
    .Z(_04644_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09667_ (.I0(_04644_),
    .I1(\soc.rom_encoder_0.request_address[2] ),
    .S(_04632_),
    .Z(_04645_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09668_ (.I(_04645_),
    .Z(_00916_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09669_ (.I(\soc.cpu.PC.REG.data[3] ),
    .ZN(_04646_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09670_ (.A1(_04639_),
    .A2(_04646_),
    .ZN(_04647_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09671_ (.A1(_04639_),
    .A2(\soc.rom_loader.current_address[3] ),
    .B(_04647_),
    .ZN(_04648_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09672_ (.A1(\soc.rom_encoder_0.request_address[3] ),
    .A2(_04618_),
    .ZN(_04649_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09673_ (.A1(_04618_),
    .A2(_04648_),
    .B(_04649_),
    .ZN(_00917_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09674_ (.I0(\soc.cpu.PC.REG.data[4] ),
    .I1(\soc.rom_loader.current_address[4] ),
    .S(_04638_),
    .Z(_04650_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09675_ (.I0(_04650_),
    .I1(\soc.rom_encoder_0.request_address[4] ),
    .S(_04632_),
    .Z(_04651_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09676_ (.I(_04651_),
    .Z(_00918_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09677_ (.I0(\soc.cpu.PC.REG.data[5] ),
    .I1(\soc.rom_loader.current_address[5] ),
    .S(_04638_),
    .Z(_04652_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09678_ (.I0(_04652_),
    .I1(\soc.rom_encoder_0.request_address[5] ),
    .S(_04632_),
    .Z(_04653_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09679_ (.I(_04653_),
    .Z(_00919_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09680_ (.A1(_04639_),
    .A2(\soc.rom_loader.current_address[6] ),
    .Z(_04654_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _09681_ (.A1(_04426_),
    .A2(\soc.cpu.PC.REG.data[6] ),
    .B(_04617_),
    .C(_04654_),
    .ZN(_04655_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09682_ (.A1(_04468_),
    .A2(_04618_),
    .B(_04655_),
    .ZN(_00920_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09683_ (.I(\soc.cpu.PC.REG.data[7] ),
    .ZN(_04656_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09684_ (.A1(_04639_),
    .A2(_04656_),
    .ZN(_04657_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09685_ (.A1(_04639_),
    .A2(\soc.rom_loader.current_address[7] ),
    .B(_04657_),
    .ZN(_04658_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09686_ (.A1(\soc.rom_encoder_0.request_address[7] ),
    .A2(_04618_),
    .ZN(_04659_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09687_ (.A1(_04618_),
    .A2(_04658_),
    .B(_04659_),
    .ZN(_00921_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09688_ (.I0(\soc.cpu.PC.REG.data[8] ),
    .I1(\soc.rom_loader.current_address[8] ),
    .S(_04638_),
    .Z(_04660_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09689_ (.I0(_04660_),
    .I1(\soc.rom_encoder_0.request_address[8] ),
    .S(_04617_),
    .Z(_04661_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09690_ (.I(_04661_),
    .Z(_00922_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09691_ (.I0(\soc.cpu.PC.REG.data[9] ),
    .I1(\soc.rom_loader.current_address[9] ),
    .S(_04638_),
    .Z(_04662_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09692_ (.I0(_04662_),
    .I1(\soc.rom_encoder_0.request_address[9] ),
    .S(_04617_),
    .Z(_04663_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09693_ (.I(_04663_),
    .Z(_00923_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09694_ (.I(\soc.cpu.PC.REG.data[10] ),
    .ZN(_04664_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09695_ (.A1(_04639_),
    .A2(_04664_),
    .ZN(_04665_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09696_ (.A1(_04639_),
    .A2(\soc.rom_loader.current_address[10] ),
    .B(_04665_),
    .ZN(_04666_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09697_ (.A1(\soc.rom_encoder_0.request_address[10] ),
    .A2(_04618_),
    .ZN(_04667_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09698_ (.A1(_04618_),
    .A2(_04666_),
    .B(_04667_),
    .ZN(_00924_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09699_ (.I0(\soc.cpu.PC.REG.data[11] ),
    .I1(\soc.rom_loader.current_address[11] ),
    .S(_04638_),
    .Z(_04668_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09700_ (.I0(_04668_),
    .I1(\soc.rom_encoder_0.request_address[11] ),
    .S(_04617_),
    .Z(_04669_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09701_ (.I(_04669_),
    .Z(_00925_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09702_ (.I0(\soc.cpu.PC.REG.data[12] ),
    .I1(\soc.rom_loader.current_address[12] ),
    .S(_04638_),
    .Z(_04670_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09703_ (.I0(_04670_),
    .I1(\soc.rom_encoder_0.request_address[12] ),
    .S(_04617_),
    .Z(_04671_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09704_ (.I(_04671_),
    .Z(_00926_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09705_ (.I0(\soc.cpu.PC.REG.data[13] ),
    .I1(\soc.rom_loader.current_address[13] ),
    .S(_04638_),
    .Z(_04672_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09706_ (.I0(_04672_),
    .I1(\soc.rom_encoder_0.request_address[13] ),
    .S(_04617_),
    .Z(_04673_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09707_ (.I(_04673_),
    .Z(_00927_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09708_ (.I0(\soc.cpu.PC.REG.data[14] ),
    .I1(\soc.rom_loader.current_address[14] ),
    .S(_04638_),
    .Z(_04674_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09709_ (.I0(_04674_),
    .I1(\soc.rom_encoder_0.request_address[14] ),
    .S(_04617_),
    .Z(_04675_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09710_ (.I(_04675_),
    .Z(_00928_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09711_ (.I(net58),
    .ZN(_04676_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _09712_ (.A1(_02548_),
    .A2(_02554_),
    .ZN(_04677_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09713_ (.A1(_02549_),
    .A2(_02553_),
    .B(_04677_),
    .ZN(_04678_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _09714_ (.A1(_02480_),
    .A2(_02481_),
    .A3(_02485_),
    .ZN(_04679_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09715_ (.A1(_02482_),
    .A2(_02499_),
    .ZN(_04680_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _09716_ (.A1(_04679_),
    .A2(_04680_),
    .A3(_03778_),
    .B(\soc.ram_encoder_0.output_buffer[16] ),
    .ZN(_04681_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09717_ (.A1(_04680_),
    .A2(_03777_),
    .B1(_03788_),
    .B2(\soc.ram_encoder_0.request_data_out[12] ),
    .ZN(_04682_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09718_ (.I(\soc.ram_encoder_0.initializing_step[2] ),
    .ZN(_04683_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09719_ (.A1(\soc.ram_encoder_0.initializing_step[1] ),
    .A2(\soc.ram_encoder_0.initializing_step[0] ),
    .ZN(_04684_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09720_ (.A1(_02548_),
    .A2(_02550_),
    .ZN(_04685_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _09721_ (.A1(_04683_),
    .A2(_02549_),
    .A3(_04684_),
    .B(_04685_),
    .ZN(_04686_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09722_ (.A1(_04681_),
    .A2(_04682_),
    .A3(_04686_),
    .ZN(_04687_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09723_ (.A1(_04678_),
    .A2(_04687_),
    .ZN(_04688_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _09724_ (.A1(_04676_),
    .A2(_04678_),
    .B(_04688_),
    .C(_01381_),
    .ZN(_00929_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _09725_ (.A1(\soc.ram_encoder_0.output_buffer[17] ),
    .A2(_03814_),
    .B1(_03788_),
    .B2(\soc.ram_encoder_0.request_data_out[13] ),
    .C(_03817_),
    .ZN(_04689_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09726_ (.A1(net59),
    .A2(_04677_),
    .ZN(_04690_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _09727_ (.A1(_04677_),
    .A2(_04689_),
    .B(_04690_),
    .C(_01381_),
    .ZN(_00930_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _09728_ (.A1(\soc.ram_encoder_0.output_buffer[18] ),
    .A2(_03814_),
    .B1(_03788_),
    .B2(\soc.ram_encoder_0.request_data_out[14] ),
    .C(_03817_),
    .ZN(_04691_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09729_ (.A1(net60),
    .A2(_04677_),
    .ZN(_04692_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _09730_ (.A1(_04677_),
    .A2(_04691_),
    .B(_04692_),
    .C(_01381_),
    .ZN(_00931_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _09731_ (.A1(\soc.ram_encoder_0.output_buffer[19] ),
    .A2(_03814_),
    .B1(_03788_),
    .B2(\soc.ram_encoder_0.request_data_out[15] ),
    .C(_03817_),
    .ZN(_04693_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09732_ (.A1(net61),
    .A2(_04677_),
    .ZN(_04694_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _09733_ (.A1(_04677_),
    .A2(_04693_),
    .B(_04694_),
    .C(_01381_),
    .ZN(_00932_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09734_ (.A1(_01445_),
    .A2(_02276_),
    .ZN(_04695_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _09735_ (.I(_04695_),
    .Z(_04696_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _09736_ (.I(_04696_),
    .Z(_04697_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09737_ (.I0(_02213_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[3][0] ),
    .S(_04697_),
    .Z(_04698_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09738_ (.I(_04698_),
    .Z(_00933_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09739_ (.I0(_02219_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[3][1] ),
    .S(_04697_),
    .Z(_04699_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09740_ (.I(_04699_),
    .Z(_00934_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09741_ (.I0(_02221_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[3][2] ),
    .S(_04697_),
    .Z(_04700_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09742_ (.I(_04700_),
    .Z(_00935_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09743_ (.I0(_02223_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[3][3] ),
    .S(_04697_),
    .Z(_04701_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09744_ (.I(_04701_),
    .Z(_00936_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09745_ (.I0(_02225_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[3][4] ),
    .S(_04697_),
    .Z(_04702_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09746_ (.I(_04702_),
    .Z(_00937_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09747_ (.I0(_02227_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[3][5] ),
    .S(_04697_),
    .Z(_04703_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09748_ (.I(_04703_),
    .Z(_00938_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09749_ (.I0(_02229_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[3][6] ),
    .S(_04697_),
    .Z(_04704_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09750_ (.I(_04704_),
    .Z(_00939_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09751_ (.I0(_02231_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[3][7] ),
    .S(_04697_),
    .Z(_04705_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09752_ (.I(_04705_),
    .Z(_00940_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09753_ (.I0(_02233_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[3][8] ),
    .S(_04697_),
    .Z(_04706_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09754_ (.I(_04706_),
    .Z(_00941_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09755_ (.I0(_02235_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[3][9] ),
    .S(_04697_),
    .Z(_04707_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09756_ (.I(_04707_),
    .Z(_00942_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _09757_ (.I(_04695_),
    .Z(_04708_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09758_ (.I0(_02237_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[3][10] ),
    .S(_04708_),
    .Z(_04709_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09759_ (.I(_04709_),
    .Z(_00943_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09760_ (.I0(_02240_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[3][11] ),
    .S(_04708_),
    .Z(_04710_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09761_ (.I(_04710_),
    .Z(_00944_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09762_ (.I0(_02242_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[3][12] ),
    .S(_04708_),
    .Z(_04711_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09763_ (.I(_04711_),
    .Z(_00945_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09764_ (.I0(_02244_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[3][13] ),
    .S(_04708_),
    .Z(_04712_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09765_ (.I(_04712_),
    .Z(_00946_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09766_ (.I0(_02246_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[3][14] ),
    .S(_04708_),
    .Z(_04713_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09767_ (.I(_04713_),
    .Z(_00947_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09768_ (.I0(_02248_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[3][15] ),
    .S(_04708_),
    .Z(_04714_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09769_ (.I(_04714_),
    .Z(_00948_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09770_ (.I0(_02250_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[3][16] ),
    .S(_04708_),
    .Z(_04715_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09771_ (.I(_04715_),
    .Z(_00949_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09772_ (.I0(_02252_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[3][17] ),
    .S(_04708_),
    .Z(_04716_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09773_ (.I(_04716_),
    .Z(_00950_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09774_ (.I0(_02254_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[3][18] ),
    .S(_04708_),
    .Z(_04717_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09775_ (.I(_04717_),
    .Z(_00951_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09776_ (.I0(_02256_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[3][19] ),
    .S(_04708_),
    .Z(_04718_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09777_ (.I(_04718_),
    .Z(_00952_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09778_ (.I0(_02258_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[3][20] ),
    .S(_04696_),
    .Z(_04719_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09779_ (.I(_04719_),
    .Z(_00953_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09780_ (.I0(_02260_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[3][21] ),
    .S(_04696_),
    .Z(_04720_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09781_ (.I(_04720_),
    .Z(_00954_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09782_ (.I0(_02262_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[3][22] ),
    .S(_04696_),
    .Z(_04721_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09783_ (.I(_04721_),
    .Z(_00955_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09784_ (.I0(_02264_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[3][23] ),
    .S(_04696_),
    .Z(_04722_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09785_ (.I(_04722_),
    .Z(_00956_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09786_ (.I0(_02266_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[3][24] ),
    .S(_04696_),
    .Z(_04723_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09787_ (.I(_04723_),
    .Z(_00957_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09788_ (.I0(_02268_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[3][25] ),
    .S(_04696_),
    .Z(_04724_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09789_ (.I(_04724_),
    .Z(_00958_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09790_ (.I0(_02270_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[3][26] ),
    .S(_04696_),
    .Z(_04725_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09791_ (.I(_04725_),
    .Z(_00959_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09792_ (.I0(_02272_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[3][27] ),
    .S(_04696_),
    .Z(_04726_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09793_ (.I(_04726_),
    .Z(_00960_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09794_ (.I0(_02274_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[3][28] ),
    .S(_04696_),
    .Z(_04727_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09795_ (.I(_04727_),
    .Z(_00961_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09796_ (.A1(\soc.rom_encoder_0.initializing_step[4] ),
    .A2(\soc.rom_encoder_0.initializing_step[2] ),
    .ZN(_04728_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09797_ (.A1(\soc.rom_encoder_0.initializing_step[3] ),
    .A2(_04728_),
    .ZN(_04729_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _09798_ (.A1(\soc.rom_encoder_0.initializing_step[1] ),
    .A2(_02459_),
    .A3(_04729_),
    .ZN(_04730_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09799_ (.A1(_02111_),
    .A2(_02456_),
    .ZN(_04731_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _09800_ (.A1(_02111_),
    .A2(_02456_),
    .A3(_02450_),
    .ZN(_04732_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09801_ (.A1(_02459_),
    .A2(_04732_),
    .ZN(_04733_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09802_ (.A1(_02459_),
    .A2(_04731_),
    .B(_04733_),
    .ZN(_04734_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09803_ (.A1(_04730_),
    .A2(_04734_),
    .B(\soc.rom_encoder_0.initialized ),
    .ZN(_04735_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09804_ (.A1(_01396_),
    .A2(_04735_),
    .ZN(_00962_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09805_ (.I(_02445_),
    .ZN(_04736_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _09806_ (.A1(_04736_),
    .A2(_02463_),
    .B1(_04566_),
    .B2(_04571_),
    .ZN(_04737_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09807_ (.A1(\soc.rom_encoder_0.toggled_sram_sck ),
    .A2(_04737_),
    .ZN(_04738_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _09808_ (.A1(_02434_),
    .A2(_02435_),
    .A3(_04738_),
    .ZN(_04739_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09809_ (.I(_04739_),
    .Z(_04740_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09810_ (.I(_04739_),
    .Z(_04741_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09811_ (.I(_04567_),
    .Z(_04742_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09812_ (.I(_04742_),
    .Z(_04743_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09813_ (.A1(\soc.rom_encoder_0.request_data_out[0] ),
    .A2(_04743_),
    .ZN(_04744_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09814_ (.A1(net5),
    .A2(_04566_),
    .ZN(_04745_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09815_ (.A1(_04741_),
    .A2(_04744_),
    .A3(_04745_),
    .ZN(_04746_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09816_ (.A1(\soc.cpu.DMuxJMP.sel[0] ),
    .A2(_04740_),
    .B(_04746_),
    .ZN(_04747_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09817_ (.A1(_01396_),
    .A2(_04747_),
    .ZN(_00963_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09818_ (.A1(\soc.rom_encoder_0.request_data_out[1] ),
    .A2(_04743_),
    .ZN(_04748_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09819_ (.A1(net6),
    .A2(_04566_),
    .ZN(_04749_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09820_ (.A1(_04741_),
    .A2(_04748_),
    .A3(_04749_),
    .ZN(_04750_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09821_ (.A1(\soc.cpu.DMuxJMP.sel[1] ),
    .A2(_04740_),
    .B(_04750_),
    .ZN(_04751_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09822_ (.A1(_01396_),
    .A2(_04751_),
    .ZN(_00964_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09823_ (.I(_01395_),
    .Z(_04752_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09824_ (.A1(\soc.rom_encoder_0.request_data_out[2] ),
    .A2(_04743_),
    .ZN(_04753_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09825_ (.A1(net7),
    .A2(_04566_),
    .ZN(_04754_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09826_ (.A1(_04741_),
    .A2(_04753_),
    .A3(_04754_),
    .ZN(_04755_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09827_ (.A1(\soc.cpu.DMuxJMP.sel[2] ),
    .A2(_04740_),
    .B(_04755_),
    .ZN(_04756_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09828_ (.A1(_04752_),
    .A2(_04756_),
    .ZN(_00965_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09829_ (.A1(\soc.rom_encoder_0.request_data_out[3] ),
    .A2(_04743_),
    .ZN(_04757_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09830_ (.A1(net8),
    .A2(_04566_),
    .ZN(_04758_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09831_ (.A1(_04741_),
    .A2(_04757_),
    .A3(_04758_),
    .ZN(_04759_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09832_ (.A1(\soc.cpu.instruction[3] ),
    .A2(_04740_),
    .B(_04759_),
    .ZN(_04760_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09833_ (.A1(_04752_),
    .A2(_04760_),
    .ZN(_00966_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09834_ (.I(_04742_),
    .Z(_04761_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09835_ (.I(_04739_),
    .Z(_04762_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09836_ (.A1(\soc.rom_encoder_0.request_data_out[4] ),
    .A2(_04743_),
    .ZN(_04763_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _09837_ (.A1(_04583_),
    .A2(_04761_),
    .B(_04762_),
    .C(_04763_),
    .ZN(_04764_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09838_ (.A1(\soc.cpu.instruction[4] ),
    .A2(_04740_),
    .B(_04764_),
    .ZN(_04765_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09839_ (.A1(_04752_),
    .A2(_04765_),
    .ZN(_00967_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09840_ (.A1(\soc.rom_encoder_0.request_data_out[5] ),
    .A2(_04743_),
    .ZN(_04766_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _09841_ (.A1(_04588_),
    .A2(_04761_),
    .B(_04762_),
    .C(_04766_),
    .ZN(_04767_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09842_ (.A1(\soc.cpu.instruction[5] ),
    .A2(_04740_),
    .B(_04767_),
    .ZN(_04768_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09843_ (.A1(_04752_),
    .A2(_04768_),
    .ZN(_00968_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09844_ (.A1(\soc.rom_encoder_0.request_data_out[6] ),
    .A2(_04743_),
    .ZN(_04769_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _09845_ (.A1(_04590_),
    .A2(_04761_),
    .B(_04762_),
    .C(_04769_),
    .ZN(_04770_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09846_ (.A1(_01615_),
    .A2(_04740_),
    .B(_04770_),
    .ZN(_04771_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09847_ (.A1(_04752_),
    .A2(_04771_),
    .ZN(_00969_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09848_ (.A1(\soc.rom_encoder_0.request_data_out[7] ),
    .A2(_04743_),
    .ZN(_04772_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _09849_ (.A1(_04592_),
    .A2(_04761_),
    .B(_04762_),
    .C(_04772_),
    .ZN(_04773_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09850_ (.A1(_01669_),
    .A2(_04740_),
    .B(_04773_),
    .ZN(_04774_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09851_ (.A1(_04752_),
    .A2(_04774_),
    .ZN(_00970_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09852_ (.A1(\soc.rom_encoder_0.request_data_out[8] ),
    .A2(_04742_),
    .ZN(_04775_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _09853_ (.A1(_04594_),
    .A2(_04761_),
    .B(_04762_),
    .C(_04775_),
    .ZN(_04776_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09854_ (.A1(_01705_),
    .A2(_04740_),
    .B(_04776_),
    .ZN(_04777_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09855_ (.A1(_04752_),
    .A2(_04777_),
    .ZN(_00971_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09856_ (.A1(\soc.rom_encoder_0.request_data_out[9] ),
    .A2(_04742_),
    .ZN(_04778_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _09857_ (.A1(_04596_),
    .A2(_04761_),
    .B(_04762_),
    .C(_04778_),
    .ZN(_04779_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09858_ (.A1(_01717_),
    .A2(_04740_),
    .B(_04779_),
    .ZN(_04780_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09859_ (.A1(_04752_),
    .A2(_04780_),
    .ZN(_00972_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09860_ (.A1(\soc.rom_encoder_0.request_data_out[10] ),
    .A2(_04742_),
    .ZN(_04781_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _09861_ (.A1(_04598_),
    .A2(_04761_),
    .B(_04762_),
    .C(_04781_),
    .ZN(_04782_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09862_ (.A1(_01702_),
    .A2(_04741_),
    .B(_04782_),
    .ZN(_04783_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09863_ (.A1(_04752_),
    .A2(_04783_),
    .ZN(_00973_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09864_ (.A1(\soc.rom_encoder_0.request_data_out[11] ),
    .A2(_04742_),
    .ZN(_04784_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _09865_ (.A1(_04600_),
    .A2(_04761_),
    .B(_04762_),
    .C(_04784_),
    .ZN(_04785_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09866_ (.A1(\soc.cpu.ALU.zx ),
    .A2(_04741_),
    .B(_04785_),
    .ZN(_04786_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09867_ (.A1(_04752_),
    .A2(_04786_),
    .ZN(_00974_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09868_ (.I(_01395_),
    .Z(_04787_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09869_ (.A1(\soc.rom_encoder_0.request_data_out[12] ),
    .A2(_04742_),
    .ZN(_04788_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _09870_ (.A1(_04603_),
    .A2(_04761_),
    .B(_04762_),
    .C(_04788_),
    .ZN(_04789_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09871_ (.A1(_01598_),
    .A2(_04741_),
    .B(_04789_),
    .ZN(_04790_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09872_ (.A1(_04787_),
    .A2(_04790_),
    .ZN(_00975_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09873_ (.A1(\soc.rom_encoder_0.request_data_out[13] ),
    .A2(_04742_),
    .ZN(_04791_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _09874_ (.A1(_04605_),
    .A2(_04761_),
    .B(_04762_),
    .C(_04791_),
    .ZN(_04792_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09875_ (.A1(\soc.cpu.instruction[13] ),
    .A2(_04741_),
    .B(_04792_),
    .ZN(_04793_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09876_ (.A1(_04787_),
    .A2(_04793_),
    .ZN(_00976_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09877_ (.A1(\soc.rom_encoder_0.request_data_out[14] ),
    .A2(_04742_),
    .ZN(_04794_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _09878_ (.A1(_04607_),
    .A2(_04743_),
    .B(_04739_),
    .C(_04794_),
    .ZN(_04795_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09879_ (.A1(\soc.cpu.instruction[14] ),
    .A2(_04741_),
    .B(_04795_),
    .ZN(_04796_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09880_ (.A1(_04787_),
    .A2(_04796_),
    .ZN(_00977_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09881_ (.A1(\soc.rom_encoder_0.request_data_out[15] ),
    .A2(_04742_),
    .ZN(_04797_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _09882_ (.A1(_04609_),
    .A2(_04743_),
    .B(_04739_),
    .C(_04797_),
    .ZN(_04798_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09883_ (.A1(_01553_),
    .A2(_04741_),
    .B(_04798_),
    .ZN(_04799_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09884_ (.A1(_04787_),
    .A2(_04799_),
    .ZN(_00978_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09885_ (.A1(_02436_),
    .A2(_02454_),
    .B(\soc.rom_encoder_0.current_state[2] ),
    .ZN(_04800_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09886_ (.A1(_04738_),
    .A2(_04800_),
    .B(net62),
    .ZN(_04801_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _09887_ (.A1(_02438_),
    .A2(_04730_),
    .B(_02450_),
    .C(_02444_),
    .ZN(_04802_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _09888_ (.A1(_04738_),
    .A2(_04800_),
    .A3(_04802_),
    .Z(_04803_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09889_ (.A1(_04254_),
    .A2(_04801_),
    .A3(_04803_),
    .ZN(_00979_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _09890_ (.A1(_02456_),
    .A2(_02448_),
    .B(_04614_),
    .C(_02443_),
    .ZN(_04804_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _09891_ (.A1(\soc.rom_encoder_0.current_state[2] ),
    .A2(_02457_),
    .A3(_04614_),
    .ZN(_04805_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09892_ (.A1(_01395_),
    .A2(_04805_),
    .ZN(_04806_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09893_ (.A1(net53),
    .A2(_04804_),
    .B(_04806_),
    .ZN(_00980_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09894_ (.A1(_02433_),
    .A2(_04730_),
    .B(_02450_),
    .ZN(_04807_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09895_ (.A1(_02437_),
    .A2(_04807_),
    .ZN(_04808_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _09896_ (.A1(_03765_),
    .A2(_04615_),
    .A3(_04737_),
    .A4(_04808_),
    .ZN(_04809_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09897_ (.A1(_04573_),
    .A2(_04809_),
    .ZN(_04810_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09898_ (.A1(_02454_),
    .A2(_04810_),
    .B(_04601_),
    .ZN(_04811_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09899_ (.A1(_02454_),
    .A2(_04810_),
    .B(_04811_),
    .ZN(_00981_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09900_ (.A1(_02436_),
    .A2(_02454_),
    .ZN(_04812_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09901_ (.A1(_04812_),
    .A2(_02525_),
    .ZN(_04813_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09902_ (.A1(_02435_),
    .A2(_04809_),
    .ZN(_04814_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _09903_ (.A1(_04809_),
    .A2(_04813_),
    .B(_04814_),
    .C(_04254_),
    .ZN(_00982_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09904_ (.A1(_04812_),
    .A2(_04809_),
    .B(\soc.rom_encoder_0.current_state[2] ),
    .ZN(_04815_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _09905_ (.A1(_02443_),
    .A2(_04809_),
    .B(_04815_),
    .C(_04254_),
    .ZN(_00983_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09906_ (.A1(_04254_),
    .A2(_04734_),
    .Z(_04816_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09907_ (.I(_04816_),
    .Z(_00984_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09908_ (.A1(_02459_),
    .A2(_04731_),
    .B(\soc.rom_encoder_0.initializing_step[1] ),
    .ZN(_04817_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09909_ (.A1(\soc.rom_encoder_0.toggled_sram_sck ),
    .A2(_02437_),
    .ZN(_04818_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09910_ (.A1(\soc.rom_encoder_0.initializing_step[1] ),
    .A2(_02459_),
    .B1(_03763_),
    .B2(_02460_),
    .ZN(_04819_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09911_ (.A1(_04818_),
    .A2(_04819_),
    .B(_04553_),
    .ZN(_04820_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09912_ (.A1(_04817_),
    .A2(_04820_),
    .ZN(_00985_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09913_ (.A1(\soc.rom_encoder_0.initializing_step[2] ),
    .A2(_04818_),
    .ZN(_04821_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09914_ (.A1(\soc.rom_encoder_0.initializing_step[2] ),
    .A2(\soc.rom_encoder_0.initializing_step[1] ),
    .A3(_02459_),
    .ZN(_04822_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09915_ (.A1(_02454_),
    .A2(_04731_),
    .A3(_04822_),
    .ZN(_04823_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09916_ (.A1(\soc.rom_encoder_0.initializing_step[1] ),
    .A2(_02459_),
    .B(\soc.rom_encoder_0.initializing_step[2] ),
    .ZN(_04824_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _09917_ (.A1(_04821_),
    .A2(_04823_),
    .B(_04824_),
    .C(_03714_),
    .ZN(_00986_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _09918_ (.A1(_02111_),
    .A2(_03763_),
    .A3(_04822_),
    .ZN(_04825_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09919_ (.A1(\soc.rom_encoder_0.initializing_step[3] ),
    .A2(_04825_),
    .ZN(_04826_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _09920_ (.A1(\soc.rom_encoder_0.initializing_step[3] ),
    .A2(\soc.rom_encoder_0.initializing_step[2] ),
    .A3(\soc.rom_encoder_0.initializing_step[1] ),
    .A4(_02459_),
    .ZN(_04827_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09921_ (.A1(_02454_),
    .A2(_04827_),
    .B(_04818_),
    .ZN(_04828_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _09922_ (.A1(_04243_),
    .A2(_04826_),
    .A3(_04828_),
    .ZN(_00987_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09923_ (.A1(\soc.rom_encoder_0.initializing_step[3] ),
    .A2(_04825_),
    .B(\soc.rom_encoder_0.initializing_step[4] ),
    .ZN(_04829_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _09924_ (.A1(\soc.rom_encoder_0.initializing_step[4] ),
    .A2(_04828_),
    .B(_04829_),
    .C(_03714_),
    .ZN(_00988_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09925_ (.A1(_04787_),
    .A2(\soc.ram_encoder_0.toggled_sram_sck ),
    .ZN(_00989_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09926_ (.A1(_02481_),
    .A2(_02482_),
    .ZN(_04830_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _09927_ (.A1(\soc.ram_encoder_0.current_state[2] ),
    .A2(_04830_),
    .ZN(_04831_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09928_ (.A1(\soc.ram_encoder_0.request_write ),
    .A2(_02503_),
    .B(_04831_),
    .ZN(_04832_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09929_ (.A1(\soc.ram_encoder_0.toggled_sram_sck ),
    .A2(_04832_),
    .ZN(_04833_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _09930_ (.A1(_02480_),
    .A2(_02498_),
    .ZN(_04834_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09931_ (.A1(\soc.ram_encoder_0.input_bits_left[3] ),
    .A2(\soc.ram_encoder_0.input_bits_left[4] ),
    .ZN(_04835_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09932_ (.A1(\soc.ram_encoder_0.input_bits_left[2] ),
    .A2(_04835_),
    .ZN(_04836_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09933_ (.A1(_04834_),
    .A2(_04836_),
    .B(_04831_),
    .ZN(_04837_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _09934_ (.A1(_01378_),
    .A2(_04833_),
    .A3(_04837_),
    .Z(_04838_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _09935_ (.A1(\soc.ram_encoder_0.input_bits_left[2] ),
    .A2(_04838_),
    .Z(_04839_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09936_ (.A1(\soc.ram_encoder_0.input_bits_left[2] ),
    .A2(_04838_),
    .ZN(_04840_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09937_ (.A1(_02480_),
    .A2(_04839_),
    .B(_04840_),
    .ZN(_00990_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _09938_ (.A1(\soc.ram_encoder_0.input_bits_left[3] ),
    .A2(_04839_),
    .Z(_04841_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _09939_ (.A1(_04834_),
    .A2(_04838_),
    .Z(_04842_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09940_ (.A1(\soc.ram_encoder_0.input_bits_left[3] ),
    .A2(_04839_),
    .ZN(_04843_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09941_ (.A1(_04841_),
    .A2(_04842_),
    .A3(_04843_),
    .ZN(_00991_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09942_ (.A1(\soc.ram_encoder_0.input_bits_left[4] ),
    .A2(_04841_),
    .ZN(_04844_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _09943_ (.A1(\soc.ram_encoder_0.input_bits_left[4] ),
    .A2(_04841_),
    .Z(_04845_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09944_ (.A1(_04842_),
    .A2(_04844_),
    .A3(_04845_),
    .ZN(_00992_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09945_ (.I(\soc.ram_encoder_0.input_buffer[0] ),
    .ZN(_04846_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _09946_ (.A1(\soc.ram_encoder_0.toggled_sram_sck ),
    .A2(_04834_),
    .ZN(_04847_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09947_ (.I(_04847_),
    .Z(_04848_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09948_ (.I(_04847_),
    .Z(_04849_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09949_ (.A1(net1),
    .A2(_04849_),
    .B(_04601_),
    .ZN(_04850_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09950_ (.A1(_04846_),
    .A2(_04848_),
    .B(_04850_),
    .ZN(_00993_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09951_ (.I(\soc.ram_encoder_0.input_buffer[1] ),
    .ZN(_04851_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09952_ (.A1(net2),
    .A2(_04849_),
    .B(_04601_),
    .ZN(_04852_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09953_ (.A1(_04851_),
    .A2(_04848_),
    .B(_04852_),
    .ZN(_00994_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09954_ (.I(\soc.ram_encoder_0.input_buffer[2] ),
    .ZN(_04853_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09955_ (.A1(net3),
    .A2(_04849_),
    .B(_04601_),
    .ZN(_04854_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09956_ (.A1(_04853_),
    .A2(_04848_),
    .B(_04854_),
    .ZN(_00995_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09957_ (.I(\soc.ram_encoder_0.input_buffer[3] ),
    .ZN(_04855_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09958_ (.A1(net4),
    .A2(_04849_),
    .B(_04601_),
    .ZN(_04856_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09959_ (.A1(_04855_),
    .A2(_04848_),
    .B(_04856_),
    .ZN(_00996_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09960_ (.I(\soc.ram_encoder_0.input_buffer[4] ),
    .ZN(_04857_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09961_ (.A1(\soc.ram_encoder_0.input_buffer[0] ),
    .A2(_04849_),
    .B(_04248_),
    .ZN(_04858_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09962_ (.A1(_04857_),
    .A2(_04848_),
    .B(_04858_),
    .ZN(_00997_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09963_ (.I(\soc.ram_encoder_0.input_buffer[5] ),
    .ZN(_04859_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09964_ (.A1(\soc.ram_encoder_0.input_buffer[1] ),
    .A2(_04849_),
    .B(_04248_),
    .ZN(_04860_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09965_ (.A1(_04859_),
    .A2(_04848_),
    .B(_04860_),
    .ZN(_00998_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09966_ (.I(\soc.ram_encoder_0.input_buffer[6] ),
    .ZN(_04861_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09967_ (.A1(\soc.ram_encoder_0.input_buffer[2] ),
    .A2(_04849_),
    .B(_04248_),
    .ZN(_04862_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09968_ (.A1(_04861_),
    .A2(_04848_),
    .B(_04862_),
    .ZN(_00999_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09969_ (.I(\soc.ram_encoder_0.input_buffer[7] ),
    .ZN(_04863_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09970_ (.A1(\soc.ram_encoder_0.input_buffer[3] ),
    .A2(_04849_),
    .B(_04248_),
    .ZN(_04864_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09971_ (.A1(_04863_),
    .A2(_04848_),
    .B(_04864_),
    .ZN(_01000_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09972_ (.I(\soc.ram_encoder_0.input_buffer[8] ),
    .ZN(_04865_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09973_ (.A1(\soc.ram_encoder_0.input_buffer[4] ),
    .A2(_04847_),
    .B(_04248_),
    .ZN(_04866_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09974_ (.A1(_04865_),
    .A2(_04848_),
    .B(_04866_),
    .ZN(_01001_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09975_ (.I(\soc.ram_encoder_0.input_buffer[9] ),
    .ZN(_04867_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09976_ (.A1(\soc.ram_encoder_0.input_buffer[5] ),
    .A2(_04847_),
    .B(_04248_),
    .ZN(_04868_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09977_ (.A1(_04867_),
    .A2(_04848_),
    .B(_04868_),
    .ZN(_01002_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09978_ (.I(\soc.ram_encoder_0.input_buffer[10] ),
    .ZN(_04869_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09979_ (.A1(\soc.ram_encoder_0.input_buffer[6] ),
    .A2(_04847_),
    .B(_04248_),
    .ZN(_04870_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09980_ (.A1(_04869_),
    .A2(_04849_),
    .B(_04870_),
    .ZN(_01003_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09981_ (.I(\soc.ram_encoder_0.input_buffer[11] ),
    .ZN(_04871_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09982_ (.A1(\soc.ram_encoder_0.input_buffer[7] ),
    .A2(_04847_),
    .B(_04248_),
    .ZN(_04872_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09983_ (.A1(_04871_),
    .A2(_04849_),
    .B(_04872_),
    .ZN(_01004_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09984_ (.A1(_02484_),
    .A2(_02486_),
    .ZN(_04873_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09985_ (.A1(_02484_),
    .A2(_02498_),
    .ZN(_04874_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09986_ (.A1(\soc.ram_step2_read_request ),
    .A2(\soc.ram_step1_write_request ),
    .B(_02053_),
    .ZN(_04875_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09987_ (.A1(_04874_),
    .A2(_04875_),
    .Z(_04876_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09988_ (.A1(_04833_),
    .A2(_04876_),
    .ZN(_04877_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _09989_ (.A1(_02504_),
    .A2(_04873_),
    .A3(_04877_),
    .ZN(_04878_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _09990_ (.A1(_04831_),
    .A2(_04878_),
    .ZN(_04879_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _09991_ (.I(_04879_),
    .Z(_04880_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09992_ (.A1(\soc.synch_hack_writeM ),
    .A2(_01579_),
    .A3(_04880_),
    .ZN(_04881_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09993_ (.A1(_03816_),
    .A2(_04880_),
    .B(_04881_),
    .ZN(_01005_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09994_ (.I0(\soc.ram_encoder_0.request_data_out[0] ),
    .I1(\soc.ram_encoder_0.data_out[0] ),
    .S(_04880_),
    .Z(_04882_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09995_ (.I(_04882_),
    .Z(_01006_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09996_ (.I0(\soc.ram_encoder_0.request_data_out[1] ),
    .I1(\soc.ram_encoder_0.data_out[1] ),
    .S(_04880_),
    .Z(_04883_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09997_ (.I(_04883_),
    .Z(_01007_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09998_ (.I0(\soc.ram_encoder_0.request_data_out[2] ),
    .I1(\soc.ram_encoder_0.data_out[2] ),
    .S(_04880_),
    .Z(_04884_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09999_ (.I(_04884_),
    .Z(_01008_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10000_ (.I0(\soc.ram_encoder_0.request_data_out[3] ),
    .I1(\soc.ram_encoder_0.data_out[3] ),
    .S(_04880_),
    .Z(_04885_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10001_ (.I(_04885_),
    .Z(_01009_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10002_ (.I0(\soc.ram_encoder_0.request_data_out[4] ),
    .I1(\soc.ram_encoder_0.data_out[4] ),
    .S(_04880_),
    .Z(_04886_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10003_ (.I(_04886_),
    .Z(_01010_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10004_ (.I0(\soc.ram_encoder_0.request_data_out[5] ),
    .I1(\soc.ram_encoder_0.data_out[5] ),
    .S(_04880_),
    .Z(_04887_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10005_ (.I(_04887_),
    .Z(_01011_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10006_ (.I0(\soc.ram_encoder_0.request_data_out[6] ),
    .I1(\soc.ram_encoder_0.data_out[6] ),
    .S(_04880_),
    .Z(_04888_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10007_ (.I(_04888_),
    .Z(_01012_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _10008_ (.I(_04879_),
    .Z(_04889_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10009_ (.I0(\soc.ram_encoder_0.request_data_out[7] ),
    .I1(\soc.ram_encoder_0.data_out[7] ),
    .S(_04889_),
    .Z(_04890_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10010_ (.I(_04890_),
    .Z(_01013_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10011_ (.I0(\soc.ram_encoder_0.request_data_out[8] ),
    .I1(\soc.ram_encoder_0.data_out[8] ),
    .S(_04889_),
    .Z(_04891_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10012_ (.I(_04891_),
    .Z(_01014_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10013_ (.I0(\soc.ram_encoder_0.request_data_out[9] ),
    .I1(\soc.ram_encoder_0.data_out[9] ),
    .S(_04889_),
    .Z(_04892_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10014_ (.I(_04892_),
    .Z(_01015_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10015_ (.I0(\soc.ram_encoder_0.request_data_out[10] ),
    .I1(\soc.ram_encoder_0.data_out[10] ),
    .S(_04889_),
    .Z(_04893_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10016_ (.I(_04893_),
    .Z(_01016_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10017_ (.I0(\soc.ram_encoder_0.request_data_out[11] ),
    .I1(\soc.ram_encoder_0.data_out[11] ),
    .S(_04889_),
    .Z(_04894_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10018_ (.I(_04894_),
    .Z(_01017_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10019_ (.I0(\soc.ram_encoder_0.request_data_out[12] ),
    .I1(\soc.ram_encoder_0.data_out[12] ),
    .S(_04889_),
    .Z(_04895_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10020_ (.I(_04895_),
    .Z(_01018_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10021_ (.I0(\soc.ram_encoder_0.request_data_out[13] ),
    .I1(\soc.ram_encoder_0.data_out[13] ),
    .S(_04889_),
    .Z(_04896_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10022_ (.I(_04896_),
    .Z(_01019_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10023_ (.I0(\soc.ram_encoder_0.request_data_out[14] ),
    .I1(\soc.ram_encoder_0.data_out[14] ),
    .S(_04889_),
    .Z(_04897_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10024_ (.I(_04897_),
    .Z(_01020_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10025_ (.I0(\soc.ram_encoder_0.request_data_out[15] ),
    .I1(\soc.ram_encoder_0.data_out[15] ),
    .S(_04889_),
    .Z(_04898_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10026_ (.I(_04898_),
    .Z(_01021_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10027_ (.I0(\soc.ram_encoder_0.request_address[0] ),
    .I1(\soc.ram_encoder_0.address[0] ),
    .S(_04889_),
    .Z(_04899_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10028_ (.I(_04899_),
    .Z(_01022_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _10029_ (.I(_04879_),
    .Z(_04900_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10030_ (.I0(\soc.ram_encoder_0.request_address[1] ),
    .I1(\soc.ram_encoder_0.address[1] ),
    .S(_04900_),
    .Z(_04901_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10031_ (.I(_04901_),
    .Z(_01023_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10032_ (.I0(\soc.ram_encoder_0.request_address[2] ),
    .I1(\soc.ram_encoder_0.address[2] ),
    .S(_04900_),
    .Z(_04902_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10033_ (.I(_04902_),
    .Z(_01024_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10034_ (.I0(\soc.ram_encoder_0.request_address[3] ),
    .I1(\soc.ram_encoder_0.address[3] ),
    .S(_04900_),
    .Z(_04903_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10035_ (.I(_04903_),
    .Z(_01025_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10036_ (.I0(\soc.ram_encoder_0.request_address[4] ),
    .I1(\soc.ram_encoder_0.address[4] ),
    .S(_04900_),
    .Z(_04904_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10037_ (.I(_04904_),
    .Z(_01026_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10038_ (.I0(\soc.ram_encoder_0.request_address[5] ),
    .I1(\soc.ram_encoder_0.address[5] ),
    .S(_04900_),
    .Z(_04905_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10039_ (.I(_04905_),
    .Z(_01027_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10040_ (.I0(\soc.ram_encoder_0.request_address[6] ),
    .I1(\soc.ram_encoder_0.address[6] ),
    .S(_04900_),
    .Z(_04906_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10041_ (.I(_04906_),
    .Z(_01028_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10042_ (.I0(\soc.ram_encoder_0.request_address[7] ),
    .I1(\soc.ram_encoder_0.address[7] ),
    .S(_04900_),
    .Z(_04907_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10043_ (.I(_04907_),
    .Z(_01029_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10044_ (.I0(\soc.ram_encoder_0.request_address[8] ),
    .I1(\soc.ram_encoder_0.address[8] ),
    .S(_04900_),
    .Z(_04908_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10045_ (.I(_04908_),
    .Z(_01030_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10046_ (.I0(\soc.ram_encoder_0.request_address[9] ),
    .I1(\soc.ram_encoder_0.address[9] ),
    .S(_04900_),
    .Z(_04909_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10047_ (.I(_04909_),
    .Z(_01031_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10048_ (.I0(\soc.ram_encoder_0.request_address[10] ),
    .I1(\soc.ram_encoder_0.address[10] ),
    .S(_04900_),
    .Z(_04910_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10049_ (.I(_04910_),
    .Z(_01032_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10050_ (.I0(\soc.ram_encoder_0.request_address[11] ),
    .I1(\soc.ram_encoder_0.address[11] ),
    .S(_04879_),
    .Z(_04911_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10051_ (.I(_04911_),
    .Z(_01033_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10052_ (.I0(\soc.ram_encoder_0.request_address[12] ),
    .I1(\soc.ram_encoder_0.address[12] ),
    .S(_04879_),
    .Z(_04912_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10053_ (.I(_04912_),
    .Z(_01034_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10054_ (.I0(\soc.ram_encoder_0.request_address[13] ),
    .I1(\soc.ram_encoder_0.address[13] ),
    .S(_04879_),
    .Z(_04913_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10055_ (.I(_04913_),
    .Z(_01035_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10056_ (.I0(\soc.ram_encoder_0.request_address[14] ),
    .I1(\soc.ram_encoder_0.address[14] ),
    .S(_04879_),
    .Z(_04914_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10057_ (.I(_04914_),
    .Z(_01036_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10058_ (.A1(\soc.ram_encoder_0.initialized ),
    .A2(_04254_),
    .ZN(_04915_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10059_ (.A1(\soc.ram_encoder_0.initializing_step[4] ),
    .A2(\soc.ram_encoder_0.initializing_step[2] ),
    .ZN(_04916_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10060_ (.A1(\soc.ram_encoder_0.initializing_step[3] ),
    .A2(_04916_),
    .A3(_04684_),
    .ZN(_04917_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10061_ (.I(_04917_),
    .ZN(_04918_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10062_ (.A1(_02112_),
    .A2(_02499_),
    .ZN(_04919_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10063_ (.I(_02550_),
    .ZN(_04920_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10064_ (.A1(_04830_),
    .A2(_04920_),
    .ZN(_04921_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10065_ (.A1(_04919_),
    .A2(_04921_),
    .B(\soc.ram_encoder_0.initializing_step[0] ),
    .ZN(_04922_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _10066_ (.A1(\soc.ram_encoder_0.initializing_step[0] ),
    .A2(_04919_),
    .B(_04922_),
    .C(_01378_),
    .ZN(_01059_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10067_ (.A1(_04918_),
    .A2(_01059_),
    .ZN(_04923_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10068_ (.A1(_04915_),
    .A2(_04923_),
    .ZN(_01037_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10069_ (.A1(_02503_),
    .A2(_04679_),
    .B1(_04834_),
    .B2(_04836_),
    .ZN(_04924_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _10070_ (.A1(\soc.ram_encoder_0.toggled_sram_sck ),
    .A2(_04924_),
    .ZN(_04925_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _10071_ (.A1(_02480_),
    .A2(_02481_),
    .A3(_04925_),
    .ZN(_04926_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10072_ (.I(_04926_),
    .Z(_04927_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10073_ (.I(_04926_),
    .Z(_04928_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _10074_ (.A1(_02484_),
    .A2(_02490_),
    .ZN(_04929_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10075_ (.I(_04929_),
    .Z(_04930_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10076_ (.A1(\soc.ram_encoder_0.request_data_out[0] ),
    .A2(_04930_),
    .ZN(_04931_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10077_ (.A1(net1),
    .A2(_04834_),
    .ZN(_04932_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10078_ (.A1(_04928_),
    .A2(_04931_),
    .A3(_04932_),
    .ZN(_04933_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10079_ (.A1(\soc.ram_data_out[0] ),
    .A2(_04927_),
    .B(_04933_),
    .ZN(_04934_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10080_ (.A1(_04787_),
    .A2(_04934_),
    .ZN(_01038_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10081_ (.A1(\soc.ram_encoder_0.request_data_out[1] ),
    .A2(_04930_),
    .ZN(_04935_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10082_ (.A1(net2),
    .A2(_04834_),
    .ZN(_04936_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10083_ (.A1(_04928_),
    .A2(_04935_),
    .A3(_04936_),
    .ZN(_04937_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10084_ (.A1(\soc.ram_data_out[1] ),
    .A2(_04927_),
    .B(_04937_),
    .ZN(_04938_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10085_ (.A1(_04787_),
    .A2(_04938_),
    .ZN(_01039_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10086_ (.A1(\soc.ram_encoder_0.request_data_out[2] ),
    .A2(_04930_),
    .ZN(_04939_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10087_ (.A1(net3),
    .A2(_04834_),
    .ZN(_04940_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10088_ (.A1(_04928_),
    .A2(_04939_),
    .A3(_04940_),
    .ZN(_04941_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10089_ (.A1(\soc.ram_data_out[2] ),
    .A2(_04927_),
    .B(_04941_),
    .ZN(_04942_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10090_ (.A1(_04787_),
    .A2(_04942_),
    .ZN(_01040_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10091_ (.A1(\soc.ram_encoder_0.request_data_out[3] ),
    .A2(_04930_),
    .ZN(_04943_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10092_ (.A1(net4),
    .A2(_04834_),
    .ZN(_04944_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10093_ (.A1(_04928_),
    .A2(_04943_),
    .A3(_04944_),
    .ZN(_04945_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10094_ (.A1(\soc.ram_data_out[3] ),
    .A2(_04927_),
    .B(_04945_),
    .ZN(_04946_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10095_ (.A1(_04787_),
    .A2(_04946_),
    .ZN(_01041_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10096_ (.I(_04929_),
    .Z(_04947_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10097_ (.I(_04926_),
    .Z(_04948_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10098_ (.A1(\soc.ram_encoder_0.request_data_out[4] ),
    .A2(_04930_),
    .ZN(_04949_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10099_ (.A1(_04846_),
    .A2(_04947_),
    .B(_04948_),
    .C(_04949_),
    .ZN(_04950_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10100_ (.A1(\soc.ram_data_out[4] ),
    .A2(_04927_),
    .B(_04950_),
    .ZN(_04951_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10101_ (.A1(_04787_),
    .A2(_04951_),
    .ZN(_01042_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10102_ (.I(_01395_),
    .Z(_04952_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10103_ (.A1(\soc.ram_encoder_0.request_data_out[5] ),
    .A2(_04930_),
    .ZN(_04953_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10104_ (.A1(_04851_),
    .A2(_04947_),
    .B(_04948_),
    .C(_04953_),
    .ZN(_04954_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10105_ (.A1(\soc.ram_data_out[5] ),
    .A2(_04927_),
    .B(_04954_),
    .ZN(_04955_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10106_ (.A1(_04952_),
    .A2(_04955_),
    .ZN(_01043_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10107_ (.A1(\soc.ram_encoder_0.request_data_out[6] ),
    .A2(_04930_),
    .ZN(_04956_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10108_ (.A1(_04853_),
    .A2(_04947_),
    .B(_04948_),
    .C(_04956_),
    .ZN(_04957_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10109_ (.A1(\soc.ram_data_out[6] ),
    .A2(_04927_),
    .B(_04957_),
    .ZN(_04958_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10110_ (.A1(_04952_),
    .A2(_04958_),
    .ZN(_01044_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10111_ (.A1(\soc.ram_encoder_0.request_data_out[7] ),
    .A2(_04930_),
    .ZN(_04959_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10112_ (.A1(_04855_),
    .A2(_04947_),
    .B(_04948_),
    .C(_04959_),
    .ZN(_04960_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10113_ (.A1(\soc.ram_data_out[7] ),
    .A2(_04927_),
    .B(_04960_),
    .ZN(_04961_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10114_ (.A1(_04952_),
    .A2(_04961_),
    .ZN(_01045_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10115_ (.A1(\soc.ram_encoder_0.request_data_out[8] ),
    .A2(_04929_),
    .ZN(_04962_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10116_ (.A1(_04857_),
    .A2(_04947_),
    .B(_04948_),
    .C(_04962_),
    .ZN(_04963_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10117_ (.A1(\soc.ram_data_out[8] ),
    .A2(_04927_),
    .B(_04963_),
    .ZN(_04964_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10118_ (.A1(_04952_),
    .A2(_04964_),
    .ZN(_01046_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10119_ (.A1(\soc.ram_encoder_0.request_data_out[9] ),
    .A2(_04929_),
    .ZN(_04965_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10120_ (.A1(_04859_),
    .A2(_04947_),
    .B(_04948_),
    .C(_04965_),
    .ZN(_04966_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10121_ (.A1(\soc.ram_data_out[9] ),
    .A2(_04927_),
    .B(_04966_),
    .ZN(_04967_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10122_ (.A1(_04952_),
    .A2(_04967_),
    .ZN(_01047_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10123_ (.A1(\soc.ram_encoder_0.request_data_out[10] ),
    .A2(_04929_),
    .ZN(_04968_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10124_ (.A1(_04861_),
    .A2(_04947_),
    .B(_04948_),
    .C(_04968_),
    .ZN(_04969_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10125_ (.A1(\soc.ram_data_out[10] ),
    .A2(_04928_),
    .B(_04969_),
    .ZN(_04970_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10126_ (.A1(_04952_),
    .A2(_04970_),
    .ZN(_01048_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10127_ (.A1(\soc.ram_encoder_0.request_data_out[11] ),
    .A2(_04929_),
    .ZN(_04971_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10128_ (.A1(_04863_),
    .A2(_04947_),
    .B(_04948_),
    .C(_04971_),
    .ZN(_04972_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10129_ (.A1(\soc.ram_data_out[11] ),
    .A2(_04928_),
    .B(_04972_),
    .ZN(_04973_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10130_ (.A1(_04952_),
    .A2(_04973_),
    .ZN(_01049_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10131_ (.A1(\soc.ram_encoder_0.request_data_out[12] ),
    .A2(_04929_),
    .ZN(_04974_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10132_ (.A1(_04865_),
    .A2(_04947_),
    .B(_04948_),
    .C(_04974_),
    .ZN(_04975_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10133_ (.A1(\soc.ram_data_out[12] ),
    .A2(_04928_),
    .B(_04975_),
    .ZN(_04976_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10134_ (.A1(_04952_),
    .A2(_04976_),
    .ZN(_01050_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10135_ (.A1(\soc.ram_encoder_0.request_data_out[13] ),
    .A2(_04929_),
    .ZN(_04977_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10136_ (.A1(_04867_),
    .A2(_04947_),
    .B(_04948_),
    .C(_04977_),
    .ZN(_04978_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10137_ (.A1(\soc.ram_data_out[13] ),
    .A2(_04928_),
    .B(_04978_),
    .ZN(_04979_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10138_ (.A1(_04952_),
    .A2(_04979_),
    .ZN(_01051_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10139_ (.A1(\soc.ram_encoder_0.request_data_out[14] ),
    .A2(_04929_),
    .ZN(_04980_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10140_ (.A1(_04869_),
    .A2(_04930_),
    .B(_04926_),
    .C(_04980_),
    .ZN(_04981_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10141_ (.A1(\soc.ram_data_out[14] ),
    .A2(_04928_),
    .B(_04981_),
    .ZN(_04982_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10142_ (.A1(_04952_),
    .A2(_04982_),
    .ZN(_01052_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10143_ (.A1(\soc.ram_encoder_0.request_data_out[15] ),
    .A2(_04929_),
    .ZN(_04983_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10144_ (.A1(_04871_),
    .A2(_04930_),
    .B(_04926_),
    .C(_04983_),
    .ZN(_04984_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10145_ (.A1(\soc.ram_data_out[15] ),
    .A2(_04928_),
    .B(_04984_),
    .ZN(_04985_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10146_ (.A1(_03714_),
    .A2(_04985_),
    .ZN(_01053_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _10147_ (.A1(_04873_),
    .A2(_04925_),
    .Z(_04986_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10148_ (.A1(_02548_),
    .A2(_04917_),
    .ZN(_04987_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _10149_ (.A1(_02484_),
    .A2(_02491_),
    .B(_02551_),
    .C(_04987_),
    .ZN(_04988_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10150_ (.A1(net81),
    .A2(_04986_),
    .B(_01395_),
    .ZN(_04989_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10151_ (.A1(_04986_),
    .A2(_04988_),
    .B(_04989_),
    .ZN(_01054_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _10152_ (.A1(\soc.ram_encoder_0.sram_sio_oe ),
    .A2(_04878_),
    .B(_04880_),
    .C(_01395_),
    .ZN(_04990_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10153_ (.I(_04990_),
    .ZN(_01055_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10154_ (.A1(_02485_),
    .A2(_04917_),
    .ZN(_04991_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _10155_ (.A1(_02499_),
    .A2(_02551_),
    .A3(_04991_),
    .ZN(_04992_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _10156_ (.A1(_03778_),
    .A2(_04876_),
    .A3(_04925_),
    .A4(_04992_),
    .ZN(_04993_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10157_ (.A1(_02504_),
    .A2(_04993_),
    .ZN(_04994_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _10158_ (.A1(\soc.ram_encoder_0.request_write ),
    .A2(_04831_),
    .B(_04874_),
    .C(_04994_),
    .ZN(_04995_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10159_ (.A1(_02482_),
    .A2(_04993_),
    .B(_04553_),
    .ZN(_04996_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10160_ (.A1(_04995_),
    .A2(_04996_),
    .ZN(_01056_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _10161_ (.A1(_02481_),
    .A2(_04993_),
    .B1(_04994_),
    .B2(_02510_),
    .ZN(_04997_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10162_ (.A1(_01381_),
    .A2(_04997_),
    .ZN(_01057_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _10163_ (.A1(_04831_),
    .A2(_04993_),
    .B1(_04994_),
    .B2(_02484_),
    .C(_01395_),
    .ZN(_04998_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10164_ (.I(_04998_),
    .ZN(_01058_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10165_ (.A1(\soc.ram_encoder_0.initializing_step[1] ),
    .A2(\soc.ram_encoder_0.initializing_step[0] ),
    .ZN(_04999_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10166_ (.A1(_02548_),
    .A2(_03777_),
    .ZN(_05000_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10167_ (.A1(_04999_),
    .A2(_05000_),
    .ZN(_05001_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10168_ (.A1(\soc.ram_encoder_0.initializing_step[0] ),
    .A2(_04919_),
    .B(\soc.ram_encoder_0.initializing_step[1] ),
    .ZN(_05002_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _10169_ (.A1(_04919_),
    .A2(_05001_),
    .B(_05002_),
    .C(_03714_),
    .ZN(_01060_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10170_ (.A1(\soc.ram_encoder_0.toggled_sram_sck ),
    .A2(_02492_),
    .ZN(_05003_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10171_ (.A1(_02485_),
    .A2(_05003_),
    .ZN(_05004_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10172_ (.A1(\soc.ram_encoder_0.initializing_step[2] ),
    .A2(\soc.ram_encoder_0.initializing_step[1] ),
    .A3(\soc.ram_encoder_0.initializing_step[0] ),
    .ZN(_05005_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10173_ (.A1(\soc.ram_encoder_0.initializing_step[2] ),
    .A2(_05003_),
    .B1(_05004_),
    .B2(_05005_),
    .ZN(_05006_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _10174_ (.A1(_04683_),
    .A2(_04999_),
    .B(_05006_),
    .C(_03714_),
    .ZN(_01061_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10175_ (.I(\soc.ram_encoder_0.initializing_step[3] ),
    .ZN(_05007_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _10176_ (.A1(_05007_),
    .A2(_05005_),
    .Z(_05008_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10177_ (.A1(\soc.ram_encoder_0.initializing_step[3] ),
    .A2(_05003_),
    .B1(_05004_),
    .B2(_05008_),
    .ZN(_05009_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _10178_ (.A1(_05007_),
    .A2(_05005_),
    .B(_05009_),
    .C(_03714_),
    .ZN(_01062_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10179_ (.A1(_05003_),
    .A2(_05008_),
    .ZN(_05010_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _10180_ (.A1(_02482_),
    .A2(_05003_),
    .B1(_05010_),
    .B2(\soc.ram_encoder_0.initializing_step[4] ),
    .C(_01380_),
    .ZN(_05011_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10181_ (.A1(\soc.ram_encoder_0.initializing_step[4] ),
    .A2(_05010_),
    .B(_05011_),
    .ZN(_01063_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10182_ (.I(\soc.hack_clock_0.counter[0] ),
    .ZN(_05012_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10183_ (.I(\soc.hack_clock_0.counter[4] ),
    .ZN(_05013_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10184_ (.A1(_05013_),
    .A2(\soc.hack_clock_0.counter[5] ),
    .ZN(_05014_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _10185_ (.A1(\soc.hack_clock_0.counter[3] ),
    .A2(\soc.hack_clock_0.counter[2] ),
    .A3(\soc.hack_clock_0.counter[6] ),
    .A4(_05014_),
    .ZN(_05015_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10186_ (.A1(\soc.hack_clock_0.counter[1] ),
    .A2(_05012_),
    .A3(_05015_),
    .ZN(_05016_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _10187_ (.A1(_01380_),
    .A2(_05016_),
    .ZN(_05017_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10188_ (.A1(\soc.hack_clock_0.counter[0] ),
    .A2(_05017_),
    .ZN(_01064_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10189_ (.A1(\soc.hack_clock_0.counter[1] ),
    .A2(\soc.hack_clock_0.counter[0] ),
    .Z(_05018_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10190_ (.A1(\soc.hack_clock_0.counter[1] ),
    .A2(\soc.hack_clock_0.counter[0] ),
    .ZN(_05019_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _10191_ (.A1(_05017_),
    .A2(_05018_),
    .A3(_05019_),
    .ZN(_01065_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10192_ (.A1(\soc.hack_clock_0.counter[2] ),
    .A2(_05018_),
    .Z(_05020_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10193_ (.A1(\soc.hack_clock_0.counter[2] ),
    .A2(_05018_),
    .ZN(_05021_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _10194_ (.A1(_05017_),
    .A2(_05020_),
    .A3(_05021_),
    .ZN(_01066_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10195_ (.A1(\soc.hack_clock_0.counter[3] ),
    .A2(_05020_),
    .Z(_05022_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10196_ (.A1(\soc.hack_clock_0.counter[3] ),
    .A2(_05020_),
    .ZN(_05023_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _10197_ (.A1(_05017_),
    .A2(_05022_),
    .A3(_05023_),
    .ZN(_01067_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10198_ (.A1(\soc.hack_clock_0.counter[4] ),
    .A2(_05022_),
    .Z(_05024_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10199_ (.A1(\soc.hack_clock_0.counter[4] ),
    .A2(_05022_),
    .ZN(_05025_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _10200_ (.A1(_05017_),
    .A2(_05024_),
    .A3(_05025_),
    .ZN(_01068_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10201_ (.A1(\soc.hack_clock_0.counter[5] ),
    .A2(_05024_),
    .ZN(_05026_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10202_ (.A1(_05017_),
    .A2(_05026_),
    .ZN(_01069_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10203_ (.A1(\soc.hack_clock_0.counter[5] ),
    .A2(_05024_),
    .ZN(_05027_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10204_ (.A1(\soc.hack_clock_0.counter[6] ),
    .A2(_05027_),
    .Z(_05028_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10205_ (.A1(_05017_),
    .A2(_05028_),
    .ZN(_01070_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _10206_ (.A1(_02179_),
    .A2(_04392_),
    .ZN(_05029_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _10207_ (.I(_05029_),
    .Z(_05030_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10208_ (.I0(_02213_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[5][0] ),
    .S(_05030_),
    .Z(_05031_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10209_ (.I(_05031_),
    .Z(_01071_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10210_ (.I0(_02219_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[5][1] ),
    .S(_05030_),
    .Z(_05032_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10211_ (.I(_05032_),
    .Z(_01072_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10212_ (.I0(_02221_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[5][2] ),
    .S(_05030_),
    .Z(_05033_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10213_ (.I(_05033_),
    .Z(_01073_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10214_ (.I0(_02223_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[5][3] ),
    .S(_05030_),
    .Z(_05034_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10215_ (.I(_05034_),
    .Z(_01074_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10216_ (.I0(_02225_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[5][4] ),
    .S(_05030_),
    .Z(_05035_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10217_ (.I(_05035_),
    .Z(_01075_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10218_ (.I0(_02227_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[5][5] ),
    .S(_05030_),
    .Z(_05036_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10219_ (.I(_05036_),
    .Z(_01076_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10220_ (.I0(_02229_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[5][6] ),
    .S(_05030_),
    .Z(_05037_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10221_ (.I(_05037_),
    .Z(_01077_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10222_ (.I0(_02231_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[5][7] ),
    .S(_05030_),
    .Z(_05038_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10223_ (.I(_05038_),
    .Z(_01078_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10224_ (.I0(_02233_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[5][8] ),
    .S(_05030_),
    .Z(_05039_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10225_ (.I(_05039_),
    .Z(_01079_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10226_ (.I0(_02235_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[5][9] ),
    .S(_05030_),
    .Z(_05040_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10227_ (.I(_05040_),
    .Z(_01080_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _10228_ (.I(_05029_),
    .Z(_05041_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10229_ (.I0(_02237_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[5][10] ),
    .S(_05041_),
    .Z(_05042_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10230_ (.I(_05042_),
    .Z(_01081_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10231_ (.I0(_02240_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[5][11] ),
    .S(_05041_),
    .Z(_05043_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10232_ (.I(_05043_),
    .Z(_01082_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10233_ (.I(_05041_),
    .Z(_05044_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10234_ (.I(_05029_),
    .Z(_05045_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10235_ (.A1(\soc.spi_video_ram_1.fifo_in_data[12] ),
    .A2(_05045_),
    .ZN(_05046_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10236_ (.A1(_03128_),
    .A2(_05044_),
    .B(_05046_),
    .ZN(_01083_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10237_ (.A1(\soc.spi_video_ram_1.fifo_in_data[13] ),
    .A2(_05045_),
    .ZN(_05047_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10238_ (.A1(_03225_),
    .A2(_05044_),
    .B(_05047_),
    .ZN(_01084_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10239_ (.A1(\soc.spi_video_ram_1.fifo_in_data[14] ),
    .A2(_05045_),
    .ZN(_05048_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10240_ (.A1(_03320_),
    .A2(_05044_),
    .B(_05048_),
    .ZN(_01085_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10241_ (.A1(\soc.spi_video_ram_1.fifo_in_data[15] ),
    .A2(_05045_),
    .ZN(_05049_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10242_ (.A1(_03419_),
    .A2(_05044_),
    .B(_05049_),
    .ZN(_01086_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10243_ (.I0(_02250_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[5][16] ),
    .S(_05041_),
    .Z(_05050_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10244_ (.I(_05050_),
    .Z(_01087_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10245_ (.I0(_02252_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[5][17] ),
    .S(_05041_),
    .Z(_05051_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10246_ (.I(_05051_),
    .Z(_01088_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10247_ (.I0(_02254_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[5][18] ),
    .S(_05041_),
    .Z(_05052_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10248_ (.I(_05052_),
    .Z(_01089_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10249_ (.I0(_02256_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[5][19] ),
    .S(_05041_),
    .Z(_05053_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10250_ (.I(_05053_),
    .Z(_01090_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10251_ (.I0(_02258_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[5][20] ),
    .S(_05041_),
    .Z(_05054_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10252_ (.I(_05054_),
    .Z(_01091_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10253_ (.A1(\soc.spi_video_ram_1.fifo_in_address[5] ),
    .A2(_05045_),
    .ZN(_05055_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10254_ (.A1(_03530_),
    .A2(_05044_),
    .B(_05055_),
    .ZN(_01092_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10255_ (.A1(\soc.spi_video_ram_1.fifo_in_address[6] ),
    .A2(_05045_),
    .ZN(_05056_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10256_ (.A1(_03504_),
    .A2(_05044_),
    .B(_05056_),
    .ZN(_01093_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10257_ (.A1(\soc.spi_video_ram_1.fifo_in_address[7] ),
    .A2(_05045_),
    .ZN(_05057_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10258_ (.A1(_03453_),
    .A2(_05044_),
    .B(_05057_),
    .ZN(_01094_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10259_ (.A1(\soc.spi_video_ram_1.fifo_in_address[8] ),
    .A2(_05045_),
    .ZN(_05058_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10260_ (.A1(_03357_),
    .A2(_05044_),
    .B(_05058_),
    .ZN(_01095_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10261_ (.A1(\soc.spi_video_ram_1.fifo_in_address[9] ),
    .A2(_05045_),
    .ZN(_05059_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10262_ (.A1(_03256_),
    .A2(_05044_),
    .B(_05059_),
    .ZN(_01096_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10263_ (.A1(\soc.spi_video_ram_1.fifo_in_address[10] ),
    .A2(_05045_),
    .ZN(_05060_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10264_ (.A1(_03178_),
    .A2(_05044_),
    .B(_05060_),
    .ZN(_01097_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10265_ (.I0(_02272_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[5][27] ),
    .S(_05041_),
    .Z(_05061_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10266_ (.I(_05061_),
    .Z(_01098_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10267_ (.I0(_02274_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[5][28] ),
    .S(_05041_),
    .Z(_05062_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10268_ (.I(_05062_),
    .Z(_01099_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10269_ (.A1(\soc.rom_encoder_0.initialized ),
    .A2(_04611_),
    .ZN(_05063_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10270_ (.A1(\soc.rom_encoder_0.write_enable ),
    .A2(net45),
    .ZN(_05064_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _10271_ (.A1(\soc.rom_loader.wait_fall_clk ),
    .A2(\soc.rom_loader.writing ),
    .A3(_05063_),
    .A4(_05064_),
    .ZN(_05065_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10272_ (.A1(\soc.rom_loader.rom_request ),
    .A2(_05065_),
    .B(_04611_),
    .ZN(_05066_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10273_ (.A1(_03714_),
    .A2(_05066_),
    .ZN(_01100_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10274_ (.A1(\soc.rom_loader.rom_request ),
    .A2(_04612_),
    .B(\soc.rom_loader.writing ),
    .ZN(_05067_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _10275_ (.A1(\soc.rom_loader.writing ),
    .A2(\soc.rom_loader.was_loading ),
    .A3(_04611_),
    .Z(_05068_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10276_ (.I(_05068_),
    .Z(_01119_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _10277_ (.A1(_04243_),
    .A2(_05067_),
    .A3(_01119_),
    .ZN(_01101_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10278_ (.A1(\soc.rom_encoder_0.toggled_sram_sck ),
    .A2(_01396_),
    .ZN(_01102_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10279_ (.A1(\soc.rom_loader.current_address[0] ),
    .A2(_01119_),
    .Z(_05069_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _10280_ (.A1(_04426_),
    .A2(\soc.rom_loader.was_loading ),
    .ZN(_05070_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10281_ (.I(_05070_),
    .Z(_05071_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10282_ (.A1(\soc.rom_loader.current_address[0] ),
    .A2(_01119_),
    .ZN(_05072_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _10283_ (.A1(_05069_),
    .A2(_05071_),
    .A3(_05072_),
    .ZN(_01103_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10284_ (.A1(\soc.rom_loader.current_address[1] ),
    .A2(_05069_),
    .B(_05070_),
    .ZN(_05073_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10285_ (.A1(\soc.rom_loader.current_address[1] ),
    .A2(_05069_),
    .B(_05073_),
    .ZN(_05074_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10286_ (.I(_05074_),
    .ZN(_01104_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10287_ (.A1(\soc.rom_loader.current_address[1] ),
    .A2(_05069_),
    .B(\soc.rom_loader.current_address[2] ),
    .ZN(_05075_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _10288_ (.A1(\soc.rom_loader.current_address[2] ),
    .A2(\soc.rom_loader.current_address[1] ),
    .A3(_05069_),
    .Z(_05076_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _10289_ (.A1(_05071_),
    .A2(_05075_),
    .A3(_05076_),
    .ZN(_01105_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10290_ (.A1(\soc.rom_loader.current_address[3] ),
    .A2(_05076_),
    .ZN(_05077_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10291_ (.A1(\soc.rom_loader.current_address[3] ),
    .A2(_05076_),
    .Z(_05078_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _10292_ (.A1(_05071_),
    .A2(_05077_),
    .A3(_05078_),
    .ZN(_01106_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10293_ (.A1(\soc.rom_loader.current_address[4] ),
    .A2(_05078_),
    .ZN(_05079_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10294_ (.A1(\soc.rom_loader.current_address[4] ),
    .A2(_05078_),
    .Z(_05080_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _10295_ (.A1(_05071_),
    .A2(_05079_),
    .A3(_05080_),
    .ZN(_01107_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10296_ (.A1(\soc.rom_loader.current_address[5] ),
    .A2(_05080_),
    .ZN(_05081_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10297_ (.A1(\soc.rom_loader.current_address[5] ),
    .A2(_05080_),
    .Z(_05082_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _10298_ (.A1(_05071_),
    .A2(_05081_),
    .A3(_05082_),
    .ZN(_01108_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10299_ (.A1(\soc.rom_loader.current_address[6] ),
    .A2(_05082_),
    .ZN(_05083_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10300_ (.A1(\soc.rom_loader.current_address[6] ),
    .A2(_05082_),
    .Z(_05084_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _10301_ (.A1(_05071_),
    .A2(_05083_),
    .A3(_05084_),
    .ZN(_01109_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10302_ (.A1(\soc.rom_loader.current_address[7] ),
    .A2(_05084_),
    .B(_05070_),
    .ZN(_05085_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10303_ (.A1(\soc.rom_loader.current_address[7] ),
    .A2(_05084_),
    .B(_05085_),
    .ZN(_05086_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10304_ (.I(_05086_),
    .ZN(_01110_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10305_ (.A1(\soc.rom_loader.current_address[7] ),
    .A2(_05084_),
    .B(\soc.rom_loader.current_address[8] ),
    .ZN(_05087_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _10306_ (.A1(\soc.rom_loader.current_address[8] ),
    .A2(\soc.rom_loader.current_address[7] ),
    .A3(_05084_),
    .Z(_05088_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _10307_ (.A1(_05071_),
    .A2(_05087_),
    .A3(_05088_),
    .ZN(_01111_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10308_ (.A1(\soc.rom_loader.current_address[9] ),
    .A2(_05088_),
    .ZN(_05089_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10309_ (.A1(\soc.rom_loader.current_address[9] ),
    .A2(_05088_),
    .Z(_05090_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _10310_ (.A1(_05071_),
    .A2(_05089_),
    .A3(_05090_),
    .ZN(_01112_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10311_ (.A1(\soc.rom_loader.current_address[10] ),
    .A2(_05090_),
    .ZN(_05091_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10312_ (.A1(\soc.rom_loader.current_address[10] ),
    .A2(_05090_),
    .Z(_05092_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _10313_ (.A1(_05071_),
    .A2(_05091_),
    .A3(_05092_),
    .ZN(_01113_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10314_ (.A1(\soc.rom_loader.current_address[11] ),
    .A2(_05092_),
    .ZN(_05093_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10315_ (.A1(\soc.rom_loader.current_address[11] ),
    .A2(_05092_),
    .Z(_05094_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _10316_ (.A1(_05070_),
    .A2(_05093_),
    .A3(_05094_),
    .ZN(_01114_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10317_ (.A1(\soc.rom_loader.current_address[12] ),
    .A2(_05094_),
    .ZN(_05095_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10318_ (.A1(\soc.rom_loader.current_address[12] ),
    .A2(_05094_),
    .Z(_05096_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _10319_ (.A1(_05070_),
    .A2(_05095_),
    .A3(_05096_),
    .ZN(_01115_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _10320_ (.A1(_04426_),
    .A2(\soc.rom_loader.was_loading ),
    .B1(_05096_),
    .B2(\soc.rom_loader.current_address[13] ),
    .ZN(_05097_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10321_ (.A1(\soc.rom_loader.current_address[13] ),
    .A2(_05096_),
    .B(_05097_),
    .ZN(_01116_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10322_ (.A1(\soc.rom_loader.current_address[13] ),
    .A2(_05096_),
    .ZN(_05098_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10323_ (.A1(\soc.rom_loader.current_address[14] ),
    .A2(_05098_),
    .Z(_05099_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10324_ (.A1(_05071_),
    .A2(_05099_),
    .ZN(_01117_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10325_ (.I(net45),
    .ZN(_05100_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10326_ (.A1(\soc.rom_loader.wait_fall_clk ),
    .A2(\soc.rom_loader.rom_request ),
    .B(_00817_),
    .ZN(_05101_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10327_ (.A1(\soc.rom_loader.wait_fall_clk ),
    .A2(_05100_),
    .B(_05101_),
    .ZN(_01118_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _10328_ (.A1(_01553_),
    .A2(\soc.cpu.instruction[4] ),
    .ZN(_05102_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10329_ (.I(_05102_),
    .Z(_05103_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10330_ (.I(_05102_),
    .Z(_05104_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10331_ (.A1(\soc.cpu.ALU.x[0] ),
    .A2(_05104_),
    .ZN(_05105_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10332_ (.A1(_01589_),
    .A2(_05103_),
    .B(_05105_),
    .ZN(_01120_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10333_ (.A1(\soc.cpu.ALU.x[1] ),
    .A2(_05104_),
    .ZN(_05106_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10334_ (.A1(_01613_),
    .A2(_05103_),
    .B(_05106_),
    .ZN(_01121_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10335_ (.A1(\soc.cpu.ALU.x[2] ),
    .A2(_05104_),
    .ZN(_05107_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10336_ (.A1(_01632_),
    .A2(_05103_),
    .B(_05107_),
    .ZN(_01122_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10337_ (.A1(\soc.cpu.ALU.x[3] ),
    .A2(_05104_),
    .ZN(_05108_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10338_ (.A1(_01652_),
    .A2(_05103_),
    .B(_05108_),
    .ZN(_01123_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10339_ (.I(_05102_),
    .Z(_05109_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10340_ (.A1(\soc.cpu.ALU.x[4] ),
    .A2(_05109_),
    .ZN(_05110_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10341_ (.A1(_01666_),
    .A2(_05103_),
    .B(_05110_),
    .ZN(_01124_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10342_ (.A1(\soc.cpu.ALU.x[5] ),
    .A2(_05109_),
    .ZN(_05111_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10343_ (.A1(_01680_),
    .A2(_05103_),
    .B(_05111_),
    .ZN(_01125_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10344_ (.A1(\soc.cpu.ALU.x[6] ),
    .A2(_05109_),
    .ZN(_05112_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10345_ (.A1(_01699_),
    .A2(_05103_),
    .B(_05112_),
    .ZN(_01126_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10346_ (.A1(\soc.cpu.ALU.x[7] ),
    .A2(_05109_),
    .ZN(_05113_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10347_ (.A1(_01713_),
    .A2(_05103_),
    .B(_05113_),
    .ZN(_01127_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10348_ (.A1(\soc.cpu.ALU.x[8] ),
    .A2(_05109_),
    .ZN(_05114_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10349_ (.A1(_01736_),
    .A2(_05103_),
    .B(_05114_),
    .ZN(_01128_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10350_ (.A1(\soc.cpu.ALU.x[9] ),
    .A2(_05109_),
    .ZN(_05115_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10351_ (.A1(_01752_),
    .A2(_05103_),
    .B(_05115_),
    .ZN(_01129_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10352_ (.A1(\soc.cpu.ALU.x[10] ),
    .A2(_05109_),
    .ZN(_05116_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10353_ (.A1(_01767_),
    .A2(_05104_),
    .B(_05116_),
    .ZN(_01130_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10354_ (.A1(\soc.cpu.ALU.x[11] ),
    .A2(_05109_),
    .ZN(_05117_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10355_ (.A1(_01779_),
    .A2(_05104_),
    .B(_05117_),
    .ZN(_01131_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10356_ (.A1(\soc.cpu.ALU.x[12] ),
    .A2(_05109_),
    .ZN(_05118_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10357_ (.A1(_01803_),
    .A2(_05104_),
    .B(_05118_),
    .ZN(_01132_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10358_ (.A1(\soc.cpu.ALU.x[13] ),
    .A2(_05109_),
    .ZN(_05119_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10359_ (.A1(_01819_),
    .A2(_05104_),
    .B(_05119_),
    .ZN(_01133_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10360_ (.A1(\soc.cpu.ALU.x[14] ),
    .A2(_05102_),
    .ZN(_05120_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10361_ (.A1(_01834_),
    .A2(_05104_),
    .B(_05120_),
    .ZN(_01134_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10362_ (.A1(\soc.cpu.ALU.x[15] ),
    .A2(_05102_),
    .ZN(_05121_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10363_ (.A1(_02539_),
    .A2(_05104_),
    .B(_05121_),
    .ZN(_01135_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10364_ (.A1(_02114_),
    .A2(_04392_),
    .ZN(_05122_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _10365_ (.I(_05122_),
    .Z(_05123_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _10366_ (.I(_05123_),
    .Z(_05124_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10367_ (.I0(_02213_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[6][0] ),
    .S(_05124_),
    .Z(_05125_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10368_ (.I(_05125_),
    .Z(_01136_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10369_ (.I0(_02219_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[6][1] ),
    .S(_05124_),
    .Z(_05126_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10370_ (.I(_05126_),
    .Z(_01137_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10371_ (.I0(_02221_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[6][2] ),
    .S(_05124_),
    .Z(_05127_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10372_ (.I(_05127_),
    .Z(_01138_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10373_ (.I0(_02223_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[6][3] ),
    .S(_05124_),
    .Z(_05128_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10374_ (.I(_05128_),
    .Z(_01139_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10375_ (.I0(_02225_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[6][4] ),
    .S(_05124_),
    .Z(_05129_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10376_ (.I(_05129_),
    .Z(_01140_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10377_ (.I0(_02227_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[6][5] ),
    .S(_05124_),
    .Z(_05130_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10378_ (.I(_05130_),
    .Z(_01141_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10379_ (.I0(_02229_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[6][6] ),
    .S(_05124_),
    .Z(_05131_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10380_ (.I(_05131_),
    .Z(_01142_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10381_ (.I0(_02231_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[6][7] ),
    .S(_05124_),
    .Z(_05132_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10382_ (.I(_05132_),
    .Z(_01143_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10383_ (.I0(_02233_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[6][8] ),
    .S(_05124_),
    .Z(_05133_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10384_ (.I(_05133_),
    .Z(_01144_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10385_ (.I0(_02235_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[6][9] ),
    .S(_05124_),
    .Z(_05134_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10386_ (.I(_05134_),
    .Z(_01145_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _10387_ (.I(_05122_),
    .Z(_05135_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10388_ (.I0(_02237_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[6][10] ),
    .S(_05135_),
    .Z(_05136_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10389_ (.I(_05136_),
    .Z(_01146_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10390_ (.I0(_02240_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[6][11] ),
    .S(_05135_),
    .Z(_05137_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10391_ (.I(_05137_),
    .Z(_01147_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10392_ (.I0(_02242_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[6][12] ),
    .S(_05135_),
    .Z(_05138_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10393_ (.I(_05138_),
    .Z(_01148_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10394_ (.I0(_02244_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[6][13] ),
    .S(_05135_),
    .Z(_05139_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10395_ (.I(_05139_),
    .Z(_01149_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10396_ (.I0(_02246_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[6][14] ),
    .S(_05135_),
    .Z(_05140_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10397_ (.I(_05140_),
    .Z(_01150_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10398_ (.I0(_02248_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[6][15] ),
    .S(_05135_),
    .Z(_05141_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10399_ (.I(_05141_),
    .Z(_01151_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10400_ (.I0(_02250_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[6][16] ),
    .S(_05135_),
    .Z(_05142_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10401_ (.I(_05142_),
    .Z(_01152_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10402_ (.I0(_02252_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[6][17] ),
    .S(_05135_),
    .Z(_05143_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10403_ (.I(_05143_),
    .Z(_01153_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10404_ (.I0(_02254_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[6][18] ),
    .S(_05135_),
    .Z(_05144_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10405_ (.I(_05144_),
    .Z(_01154_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10406_ (.I0(_02256_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[6][19] ),
    .S(_05135_),
    .Z(_05145_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10407_ (.I(_05145_),
    .Z(_01155_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10408_ (.I0(_02258_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[6][20] ),
    .S(_05123_),
    .Z(_05146_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10409_ (.I(_05146_),
    .Z(_01156_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10410_ (.I0(_02260_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[6][21] ),
    .S(_05123_),
    .Z(_05147_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10411_ (.I(_05147_),
    .Z(_01157_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10412_ (.I0(_02262_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[6][22] ),
    .S(_05123_),
    .Z(_05148_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10413_ (.I(_05148_),
    .Z(_01158_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10414_ (.I0(_02264_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[6][23] ),
    .S(_05123_),
    .Z(_05149_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10415_ (.I(_05149_),
    .Z(_01159_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10416_ (.I0(_02266_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[6][24] ),
    .S(_05123_),
    .Z(_05150_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10417_ (.I(_05150_),
    .Z(_01160_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10418_ (.I0(_02268_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[6][25] ),
    .S(_05123_),
    .Z(_05151_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10419_ (.I(_05151_),
    .Z(_01161_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10420_ (.I0(_02270_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[6][26] ),
    .S(_05123_),
    .Z(_05152_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10421_ (.I(_05152_),
    .Z(_01162_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10422_ (.I0(_02272_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[6][27] ),
    .S(_05123_),
    .Z(_05153_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10423_ (.I(_05153_),
    .Z(_01163_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10424_ (.I0(_02274_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[6][28] ),
    .S(_05123_),
    .Z(_05154_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10425_ (.I(_05154_),
    .Z(_01164_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10426_ (.A1(_01378_),
    .A2(_05016_),
    .ZN(_05155_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10427_ (.I(_05155_),
    .Z(_01181_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10428_ (.A1(net90),
    .A2(_01181_),
    .ZN(_05156_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10429_ (.A1(net90),
    .A2(_05017_),
    .B(_05156_),
    .ZN(_01165_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10430_ (.A1(_01615_),
    .A2(_01751_),
    .Z(_05157_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10431_ (.A1(_01615_),
    .A2(_01766_),
    .Z(_05158_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10432_ (.A1(_01615_),
    .A2(_01802_),
    .Z(_05159_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _10433_ (.A1(_01589_),
    .A2(_01613_),
    .A3(_01632_),
    .A4(_01652_),
    .Z(_05160_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _10434_ (.A1(_01666_),
    .A2(_01680_),
    .A3(_01713_),
    .A4(_05160_),
    .Z(_05161_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10435_ (.A1(_01699_),
    .A2(_01736_),
    .A3(_05161_),
    .ZN(_05162_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _10436_ (.A1(_05157_),
    .A2(_05158_),
    .A3(_05159_),
    .A4(_05162_),
    .ZN(_05163_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _10437_ (.A1(_01779_),
    .A2(_01819_),
    .A3(_05163_),
    .Z(_05164_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _10438_ (.A1(_01834_),
    .A2(_05164_),
    .B(_01554_),
    .ZN(_05165_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10439_ (.I(\soc.cpu.DMuxJMP.sel[1] ),
    .ZN(_05166_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10440_ (.A1(_01615_),
    .A2(_01833_),
    .Z(_05167_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10441_ (.A1(_01779_),
    .A2(_01819_),
    .A3(_05163_),
    .ZN(_05168_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _10442_ (.A1(_05166_),
    .A2(_05167_),
    .A3(_05168_),
    .B(_02539_),
    .ZN(_05169_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_4 _10443_ (.A1(\soc.cpu.DMuxJMP.sel[2] ),
    .A2(_02539_),
    .B1(_05165_),
    .B2(_05169_),
    .C(_01552_),
    .ZN(_05170_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10444_ (.I(_05170_),
    .Z(_05171_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10445_ (.I(_05170_),
    .Z(_05172_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10446_ (.I(_02053_),
    .Z(_05173_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10447_ (.A1(\soc.cpu.PC.in[0] ),
    .A2(_05172_),
    .B(_05173_),
    .ZN(_05174_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10448_ (.A1(\soc.cpu.PC.REG.data[0] ),
    .A2(_05171_),
    .B(_05174_),
    .ZN(_01166_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10449_ (.A1(\soc.cpu.PC.REG.data[0] ),
    .A2(\soc.cpu.PC.REG.data[1] ),
    .ZN(_05175_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10450_ (.A1(\soc.cpu.PC.in[1] ),
    .A2(_05172_),
    .B(_05173_),
    .ZN(_05176_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10451_ (.A1(_05171_),
    .A2(_05175_),
    .B(_05176_),
    .ZN(_01167_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10452_ (.A1(\soc.cpu.PC.REG.data[0] ),
    .A2(\soc.cpu.PC.REG.data[1] ),
    .ZN(_05177_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10453_ (.A1(\soc.cpu.PC.REG.data[2] ),
    .A2(_05177_),
    .Z(_05178_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10454_ (.A1(\soc.cpu.PC.in[2] ),
    .A2(_05172_),
    .B(_05173_),
    .ZN(_05179_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10455_ (.A1(_05171_),
    .A2(_05178_),
    .B(_05179_),
    .ZN(_01168_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10456_ (.A1(\soc.cpu.PC.REG.data[0] ),
    .A2(\soc.cpu.PC.REG.data[1] ),
    .A3(\soc.cpu.PC.REG.data[2] ),
    .ZN(_05180_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10457_ (.A1(\soc.cpu.PC.REG.data[3] ),
    .A2(_05180_),
    .Z(_05181_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10458_ (.A1(\soc.cpu.PC.in[3] ),
    .A2(_05172_),
    .B(_05173_),
    .ZN(_05182_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10459_ (.A1(_05171_),
    .A2(_05181_),
    .B(_05182_),
    .ZN(_01169_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10460_ (.A1(_04646_),
    .A2(_05180_),
    .ZN(_05183_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10461_ (.A1(\soc.cpu.PC.REG.data[4] ),
    .A2(_05183_),
    .ZN(_05184_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10462_ (.A1(\soc.cpu.PC.in[4] ),
    .A2(_05172_),
    .B(_05173_),
    .ZN(_05185_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10463_ (.A1(_05171_),
    .A2(_05184_),
    .B(_05185_),
    .ZN(_01170_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10464_ (.A1(\soc.cpu.PC.REG.data[4] ),
    .A2(_05183_),
    .Z(_05186_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10465_ (.A1(\soc.cpu.PC.REG.data[5] ),
    .A2(_05186_),
    .ZN(_05187_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10466_ (.I(_05170_),
    .Z(_05188_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10467_ (.A1(\soc.cpu.PC.in[5] ),
    .A2(_05188_),
    .B(_05173_),
    .ZN(_05189_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10468_ (.A1(_05171_),
    .A2(_05187_),
    .B(_05189_),
    .ZN(_01171_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10469_ (.A1(\soc.cpu.PC.REG.data[5] ),
    .A2(_05186_),
    .ZN(_05190_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10470_ (.A1(\soc.cpu.PC.REG.data[6] ),
    .A2(_05190_),
    .Z(_05191_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10471_ (.A1(\soc.cpu.PC.in[6] ),
    .A2(_05188_),
    .B(_05173_),
    .ZN(_05192_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10472_ (.A1(_05171_),
    .A2(_05191_),
    .B(_05192_),
    .ZN(_01172_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10473_ (.A1(\soc.cpu.PC.REG.data[5] ),
    .A2(\soc.cpu.PC.REG.data[6] ),
    .A3(_05186_),
    .ZN(_05193_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10474_ (.A1(\soc.cpu.PC.REG.data[7] ),
    .A2(_05193_),
    .Z(_05194_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10475_ (.A1(\soc.cpu.PC.in[7] ),
    .A2(_05188_),
    .B(_05173_),
    .ZN(_05195_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10476_ (.A1(_05171_),
    .A2(_05194_),
    .B(_05195_),
    .ZN(_01173_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10477_ (.A1(_04656_),
    .A2(_05193_),
    .ZN(_05196_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10478_ (.A1(\soc.cpu.PC.REG.data[8] ),
    .A2(_05196_),
    .ZN(_05197_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10479_ (.A1(\soc.cpu.PC.in[8] ),
    .A2(_05188_),
    .B(_05173_),
    .ZN(_05198_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10480_ (.A1(_05171_),
    .A2(_05197_),
    .B(_05198_),
    .ZN(_01174_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10481_ (.A1(\soc.cpu.PC.REG.data[8] ),
    .A2(_05196_),
    .ZN(_05199_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10482_ (.A1(\soc.cpu.PC.REG.data[9] ),
    .A2(_05199_),
    .Z(_05200_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10483_ (.I(_02053_),
    .Z(_05201_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10484_ (.A1(\soc.cpu.PC.in[9] ),
    .A2(_05188_),
    .B(_05201_),
    .ZN(_05202_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10485_ (.A1(_05171_),
    .A2(_05200_),
    .B(_05202_),
    .ZN(_01175_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10486_ (.A1(\soc.cpu.PC.REG.data[8] ),
    .A2(\soc.cpu.PC.REG.data[9] ),
    .A3(_05196_),
    .ZN(_05203_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10487_ (.A1(\soc.cpu.PC.REG.data[10] ),
    .A2(_05203_),
    .Z(_05204_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10488_ (.A1(\soc.cpu.PC.in[10] ),
    .A2(_05188_),
    .B(_05201_),
    .ZN(_05205_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10489_ (.A1(_05172_),
    .A2(_05204_),
    .B(_05205_),
    .ZN(_01176_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _10490_ (.A1(_04664_),
    .A2(_05203_),
    .ZN(_05206_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10491_ (.A1(\soc.cpu.PC.REG.data[11] ),
    .A2(_05206_),
    .ZN(_05207_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10492_ (.A1(\soc.cpu.PC.in[11] ),
    .A2(_05188_),
    .B(_05201_),
    .ZN(_05208_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10493_ (.A1(_05172_),
    .A2(_05207_),
    .B(_05208_),
    .ZN(_01177_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10494_ (.A1(\soc.cpu.PC.REG.data[11] ),
    .A2(_05206_),
    .ZN(_05209_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10495_ (.A1(\soc.cpu.PC.REG.data[12] ),
    .A2(_05209_),
    .Z(_05210_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10496_ (.A1(\soc.cpu.PC.in[12] ),
    .A2(_05188_),
    .B(_05201_),
    .ZN(_05211_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10497_ (.A1(_05172_),
    .A2(_05210_),
    .B(_05211_),
    .ZN(_01178_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10498_ (.A1(\soc.cpu.PC.REG.data[11] ),
    .A2(\soc.cpu.PC.REG.data[12] ),
    .A3(_05206_),
    .ZN(_05212_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10499_ (.A1(\soc.cpu.PC.REG.data[13] ),
    .A2(_05212_),
    .Z(_05213_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10500_ (.A1(\soc.cpu.PC.in[13] ),
    .A2(_05188_),
    .B(_05201_),
    .ZN(_05214_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10501_ (.A1(_05172_),
    .A2(_05213_),
    .B(_05214_),
    .ZN(_01179_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _10502_ (.A1(\soc.cpu.PC.REG.data[11] ),
    .A2(\soc.cpu.PC.REG.data[12] ),
    .A3(\soc.cpu.PC.REG.data[13] ),
    .A4(_05206_),
    .ZN(_05215_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10503_ (.A1(\soc.cpu.PC.REG.data[14] ),
    .A2(_05215_),
    .Z(_05216_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10504_ (.A1(\soc.cpu.PC.in[14] ),
    .A2(_05188_),
    .B(_05201_),
    .ZN(_05217_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10505_ (.A1(_05172_),
    .A2(_05216_),
    .B(_05217_),
    .ZN(_01180_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10506_ (.I(net90),
    .ZN(_05218_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10507_ (.A1(_05218_),
    .A2(_05015_),
    .A3(_05019_),
    .ZN(_05219_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _10508_ (.A1(_01455_),
    .A2(_05219_),
    .Z(_05220_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10509_ (.I(_05220_),
    .Z(_05221_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10510_ (.I(_05221_),
    .Z(_05222_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10511_ (.A1(_05015_),
    .A2(_05019_),
    .ZN(_05223_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10512_ (.A1(_05218_),
    .A2(\soc.hack_clk_strobe ),
    .A3(_05223_),
    .ZN(_05224_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10513_ (.A1(\soc.synch_hack_writeM ),
    .A2(_05224_),
    .ZN(_05225_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10514_ (.A1(_05222_),
    .A2(_05225_),
    .ZN(_01182_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10515_ (.A1(_05221_),
    .A2(_05224_),
    .ZN(_05226_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _10516_ (.I(_05226_),
    .Z(_05227_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10517_ (.I(_05227_),
    .Z(_05228_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10518_ (.A1(\soc.ram_encoder_0.address[0] ),
    .A2(_05228_),
    .ZN(_05229_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10519_ (.A1(_01564_),
    .A2(_05228_),
    .B(_05229_),
    .ZN(_01183_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10520_ (.A1(\soc.ram_encoder_0.address[1] ),
    .A2(_05228_),
    .ZN(_05230_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10521_ (.A1(_01565_),
    .A2(_05228_),
    .B(_05230_),
    .ZN(_01184_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10522_ (.A1(\soc.ram_encoder_0.address[2] ),
    .A2(_05228_),
    .ZN(_05231_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10523_ (.A1(_01619_),
    .A2(_05228_),
    .B(_05231_),
    .ZN(_01185_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10524_ (.I0(\soc.ram_encoder_0.address[3] ),
    .I1(\soc.cpu.AReg.data[3] ),
    .S(_05228_),
    .Z(_05232_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10525_ (.I(_05232_),
    .Z(_01186_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10526_ (.I0(\soc.ram_encoder_0.address[4] ),
    .I1(\soc.cpu.AReg.data[4] ),
    .S(_05228_),
    .Z(_05233_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10527_ (.I(_05233_),
    .Z(_01187_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10528_ (.I0(\soc.ram_encoder_0.address[5] ),
    .I1(\soc.cpu.AReg.data[5] ),
    .S(_05227_),
    .Z(_05234_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10529_ (.I(_05234_),
    .Z(_01188_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10530_ (.I0(\soc.ram_encoder_0.address[6] ),
    .I1(\soc.cpu.AReg.data[6] ),
    .S(_05227_),
    .Z(_05235_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10531_ (.I(_05235_),
    .Z(_01189_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10532_ (.I0(\soc.ram_encoder_0.address[7] ),
    .I1(\soc.cpu.AReg.data[7] ),
    .S(_05227_),
    .Z(_05236_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10533_ (.I(_05236_),
    .Z(_01190_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10534_ (.I0(\soc.ram_encoder_0.address[8] ),
    .I1(\soc.cpu.AReg.data[8] ),
    .S(_05227_),
    .Z(_05237_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10535_ (.I(_05237_),
    .Z(_01191_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10536_ (.I0(\soc.ram_encoder_0.address[9] ),
    .I1(\soc.cpu.AReg.data[9] ),
    .S(_05227_),
    .Z(_05238_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10537_ (.I(_05238_),
    .Z(_01192_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10538_ (.I0(\soc.ram_encoder_0.address[10] ),
    .I1(\soc.cpu.AReg.data[10] ),
    .S(_05227_),
    .Z(_05239_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10539_ (.I(_05239_),
    .Z(_01193_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10540_ (.I0(\soc.ram_encoder_0.address[11] ),
    .I1(\soc.cpu.AReg.data[11] ),
    .S(_05227_),
    .Z(_05240_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10541_ (.I(_05240_),
    .Z(_01194_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10542_ (.I0(\soc.ram_encoder_0.address[12] ),
    .I1(\soc.cpu.AReg.data[12] ),
    .S(_05227_),
    .Z(_05241_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10543_ (.I(_05241_),
    .Z(_01195_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10544_ (.A1(\soc.ram_encoder_0.address[13] ),
    .A2(_05228_),
    .ZN(_05242_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10545_ (.A1(_01456_),
    .A2(_05228_),
    .B(_05242_),
    .ZN(_01196_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10546_ (.I0(\soc.ram_encoder_0.address[14] ),
    .I1(\soc.cpu.AReg.data[14] ),
    .S(_05227_),
    .Z(_05243_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10547_ (.I(_05243_),
    .Z(_01197_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10548_ (.I(_05224_),
    .ZN(_01198_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10549_ (.I(_05222_),
    .ZN(_01199_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10550_ (.A1(_05218_),
    .A2(\soc.hack_clk_strobe ),
    .ZN(_05244_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10551_ (.A1(_05063_),
    .A2(_05244_),
    .ZN(_01200_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10552_ (.A1(_04639_),
    .A2(net45),
    .B(\soc.boot_loading_offset[0] ),
    .ZN(_05245_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _10553_ (.A1(_01895_),
    .A2(_05064_),
    .ZN(_05246_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _10554_ (.A1(_04243_),
    .A2(_05245_),
    .A3(_05246_),
    .ZN(_01201_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10555_ (.A1(\soc.boot_loading_offset[1] ),
    .A2(_05246_),
    .B(_01395_),
    .ZN(_05247_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10556_ (.A1(\soc.boot_loading_offset[1] ),
    .A2(_05246_),
    .B(_05247_),
    .ZN(_05248_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10557_ (.I(_05248_),
    .ZN(_01202_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10558_ (.A1(\soc.boot_loading_offset[1] ),
    .A2(_05246_),
    .B(\soc.boot_loading_offset[2] ),
    .ZN(_05249_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _10559_ (.A1(\soc.boot_loading_offset[2] ),
    .A2(\soc.boot_loading_offset[1] ),
    .A3(_05246_),
    .Z(_05250_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _10560_ (.A1(_04243_),
    .A2(_05249_),
    .A3(_05250_),
    .ZN(_01203_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10561_ (.A1(\soc.boot_loading_offset[3] ),
    .A2(_05250_),
    .B(_04248_),
    .ZN(_05251_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10562_ (.A1(\soc.boot_loading_offset[3] ),
    .A2(_05250_),
    .B(_05251_),
    .ZN(_01204_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10563_ (.A1(\soc.boot_loading_offset[3] ),
    .A2(_05250_),
    .ZN(_05252_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10564_ (.A1(\soc.boot_loading_offset[4] ),
    .A2(_05252_),
    .Z(_05253_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10565_ (.A1(_03714_),
    .A2(_05253_),
    .ZN(_01205_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10566_ (.A1(net90),
    .A2(\soc.hack_clk_strobe ),
    .ZN(_05254_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10567_ (.I(net19),
    .ZN(_05255_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10568_ (.A1(_05173_),
    .A2(_05254_),
    .B(_05255_),
    .ZN(_01206_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10569_ (.A1(\soc.hack_wait_clocks[0] ),
    .A2(_05254_),
    .ZN(_05256_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10570_ (.A1(\soc.hack_wait_clocks[0] ),
    .A2(_05254_),
    .ZN(_05257_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10571_ (.A1(\soc.hack_wait_clocks[1] ),
    .A2(_05257_),
    .ZN(_05258_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10572_ (.A1(_05256_),
    .A2(_05258_),
    .B(_01452_),
    .ZN(_01207_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10573_ (.I(\soc.hack_wait_clocks[1] ),
    .ZN(_05259_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10574_ (.I(_01452_),
    .ZN(_05260_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10575_ (.A1(_05259_),
    .A2(_05257_),
    .B(_05260_),
    .ZN(_01208_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _10576_ (.A1(\soc.cpu.AReg.data[0] ),
    .A2(_01455_),
    .A3(_01572_),
    .A4(_01641_),
    .ZN(_05261_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10577_ (.A1(net77),
    .A2(_05261_),
    .B(_05201_),
    .ZN(_05262_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10578_ (.A1(_01589_),
    .A2(_05261_),
    .B(_05262_),
    .ZN(_01209_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10579_ (.A1(net78),
    .A2(_05261_),
    .B(_05201_),
    .ZN(_05263_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10580_ (.A1(_01613_),
    .A2(_05261_),
    .B(_05263_),
    .ZN(_01210_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10581_ (.A1(net79),
    .A2(_05261_),
    .B(_05201_),
    .ZN(_05264_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10582_ (.A1(_01632_),
    .A2(_05261_),
    .B(_05264_),
    .ZN(_01211_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10583_ (.A1(net80),
    .A2(_05261_),
    .B(_05201_),
    .ZN(_05265_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10584_ (.A1(_01652_),
    .A2(_05261_),
    .B(_05265_),
    .ZN(_01212_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10585_ (.I(net14),
    .ZN(_05266_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10586_ (.A1(_01455_),
    .A2(_01575_),
    .Z(_05267_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10587_ (.I(_05267_),
    .Z(_05268_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10588_ (.A1(\soc.gpio_i_stored[0] ),
    .A2(_05268_),
    .B(_02053_),
    .ZN(_05269_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10589_ (.A1(_05266_),
    .A2(_05268_),
    .B(_05269_),
    .ZN(_01213_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10590_ (.I(net15),
    .ZN(_05270_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10591_ (.A1(\soc.gpio_i_stored[1] ),
    .A2(_05268_),
    .B(_02053_),
    .ZN(_05271_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10592_ (.A1(_05270_),
    .A2(_05268_),
    .B(_05271_),
    .ZN(_01214_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10593_ (.I(net16),
    .ZN(_05272_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10594_ (.A1(\soc.gpio_i_stored[2] ),
    .A2(_05268_),
    .B(_02053_),
    .ZN(_05273_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10595_ (.A1(_05272_),
    .A2(_05268_),
    .B(_05273_),
    .ZN(_01215_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10596_ (.I(net17),
    .ZN(_05274_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10597_ (.A1(\soc.gpio_i_stored[3] ),
    .A2(_05268_),
    .B(_02053_),
    .ZN(_05275_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10598_ (.A1(_05274_),
    .A2(_05268_),
    .B(_05275_),
    .ZN(_01216_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10599_ (.A1(_01445_),
    .A2(_02117_),
    .Z(_05276_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _10600_ (.I(_05276_),
    .Z(_05277_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _10601_ (.I(_05277_),
    .Z(_05278_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10602_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[19][0] ),
    .I1(\soc.spi_video_ram_1.fifo_in_data[0] ),
    .S(_05278_),
    .Z(_05279_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10603_ (.I(_05279_),
    .Z(_01217_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10604_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[19][1] ),
    .I1(_02393_),
    .S(_05278_),
    .Z(_05280_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10605_ (.I(_05280_),
    .Z(_01218_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10606_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[19][2] ),
    .I1(_02395_),
    .S(_05278_),
    .Z(_05281_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10607_ (.I(_05281_),
    .Z(_01219_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10608_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[19][3] ),
    .I1(_02397_),
    .S(_05278_),
    .Z(_05282_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10609_ (.I(_05282_),
    .Z(_01220_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10610_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[19][4] ),
    .I1(_02399_),
    .S(_05278_),
    .Z(_05283_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10611_ (.I(_05283_),
    .Z(_01221_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10612_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[19][5] ),
    .I1(_02401_),
    .S(_05278_),
    .Z(_05284_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10613_ (.I(_05284_),
    .Z(_01222_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10614_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[19][6] ),
    .I1(_02403_),
    .S(_05278_),
    .Z(_05285_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10615_ (.I(_05285_),
    .Z(_01223_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10616_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[19][7] ),
    .I1(_02405_),
    .S(_05278_),
    .Z(_05286_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10617_ (.I(_05286_),
    .Z(_01224_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10618_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[19][8] ),
    .I1(_02407_),
    .S(_05278_),
    .Z(_05287_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10619_ (.I(_05287_),
    .Z(_01225_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10620_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[19][9] ),
    .I1(_02409_),
    .S(_05278_),
    .Z(_05288_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10621_ (.I(_05288_),
    .Z(_01226_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _10622_ (.I(_05276_),
    .Z(_05289_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10623_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[19][10] ),
    .I1(_02411_),
    .S(_05289_),
    .Z(_05290_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10624_ (.I(_05290_),
    .Z(_01227_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10625_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[19][11] ),
    .I1(_02414_),
    .S(_05289_),
    .Z(_05291_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10626_ (.I(_05291_),
    .Z(_01228_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10627_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[19][12] ),
    .I1(_04047_),
    .S(_05289_),
    .Z(_05292_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10628_ (.I(_05292_),
    .Z(_01229_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10629_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[19][13] ),
    .I1(_04050_),
    .S(_05289_),
    .Z(_05293_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10630_ (.I(_05293_),
    .Z(_01230_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10631_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[19][14] ),
    .I1(_04052_),
    .S(_05289_),
    .Z(_05294_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10632_ (.I(_05294_),
    .Z(_01231_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10633_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[19][15] ),
    .I1(_04054_),
    .S(_05289_),
    .Z(_05295_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10634_ (.I(_05295_),
    .Z(_01232_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10635_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[19][16] ),
    .I1(\soc.spi_video_ram_1.fifo_in_address[0] ),
    .S(_05289_),
    .Z(_05296_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10636_ (.I(_05296_),
    .Z(_01233_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10637_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[19][17] ),
    .I1(\soc.spi_video_ram_1.fifo_in_address[1] ),
    .S(_05289_),
    .Z(_05297_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10638_ (.I(_05297_),
    .Z(_01234_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10639_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[19][18] ),
    .I1(\soc.spi_video_ram_1.fifo_in_address[2] ),
    .S(_05289_),
    .Z(_05298_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10640_ (.I(_05298_),
    .Z(_01235_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10641_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[19][19] ),
    .I1(\soc.spi_video_ram_1.fifo_in_address[3] ),
    .S(_05289_),
    .Z(_05299_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10642_ (.I(_05299_),
    .Z(_01236_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10643_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[19][20] ),
    .I1(\soc.spi_video_ram_1.fifo_in_address[4] ),
    .S(_05277_),
    .Z(_05300_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10644_ (.I(_05300_),
    .Z(_01237_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10645_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[19][21] ),
    .I1(_04061_),
    .S(_05277_),
    .Z(_05301_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10646_ (.I(_05301_),
    .Z(_01238_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10647_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[19][22] ),
    .I1(_04063_),
    .S(_05277_),
    .Z(_05302_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10648_ (.I(_05302_),
    .Z(_01239_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10649_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[19][23] ),
    .I1(_04065_),
    .S(_05277_),
    .Z(_05303_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10650_ (.I(_05303_),
    .Z(_01240_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10651_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[19][24] ),
    .I1(_04067_),
    .S(_05277_),
    .Z(_05304_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10652_ (.I(_05304_),
    .Z(_01241_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10653_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[19][25] ),
    .I1(_04069_),
    .S(_05277_),
    .Z(_05305_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10654_ (.I(_05305_),
    .Z(_01242_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10655_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[19][26] ),
    .I1(_03927_),
    .S(_05277_),
    .Z(_05306_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10656_ (.I(_05306_),
    .Z(_01243_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10657_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[19][27] ),
    .I1(\soc.spi_video_ram_1.fifo_in_address[11] ),
    .S(_05277_),
    .Z(_05307_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10658_ (.I(_05307_),
    .Z(_01244_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10659_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[19][28] ),
    .I1(\soc.spi_video_ram_1.fifo_in_address[12] ),
    .S(_05277_),
    .Z(_05308_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10660_ (.I(_05308_),
    .Z(_01245_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10661_ (.A1(_03931_),
    .A2(_02179_),
    .ZN(_05309_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _10662_ (.I(_05309_),
    .Z(_05310_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10663_ (.I0(_02213_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[29][0] ),
    .S(_05310_),
    .Z(_05311_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10664_ (.I(_05311_),
    .Z(_01246_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10665_ (.I0(_02219_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[29][1] ),
    .S(_05310_),
    .Z(_05312_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10666_ (.I(_05312_),
    .Z(_01247_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10667_ (.I0(_02221_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[29][2] ),
    .S(_05310_),
    .Z(_05313_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10668_ (.I(_05313_),
    .Z(_01248_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10669_ (.I0(_02223_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[29][3] ),
    .S(_05310_),
    .Z(_05314_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10670_ (.I(_05314_),
    .Z(_01249_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10671_ (.I0(_02225_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[29][4] ),
    .S(_05310_),
    .Z(_05315_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10672_ (.I(_05315_),
    .Z(_01250_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10673_ (.I0(_02227_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[29][5] ),
    .S(_05310_),
    .Z(_05316_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10674_ (.I(_05316_),
    .Z(_01251_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10675_ (.I0(_02229_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[29][6] ),
    .S(_05310_),
    .Z(_05317_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10676_ (.I(_05317_),
    .Z(_01252_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10677_ (.I0(_02231_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[29][7] ),
    .S(_05310_),
    .Z(_05318_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10678_ (.I(_05318_),
    .Z(_01253_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10679_ (.I0(_02233_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[29][8] ),
    .S(_05310_),
    .Z(_05319_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10680_ (.I(_05319_),
    .Z(_01254_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10681_ (.I0(_02235_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[29][9] ),
    .S(_05310_),
    .Z(_05320_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10682_ (.I(_05320_),
    .Z(_01255_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _10683_ (.I(_05309_),
    .Z(_05321_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10684_ (.I0(_02237_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[29][10] ),
    .S(_05321_),
    .Z(_05322_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10685_ (.I(_05322_),
    .Z(_01256_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10686_ (.I0(_02240_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[29][11] ),
    .S(_05321_),
    .Z(_05323_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10687_ (.I(_05323_),
    .Z(_01257_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10688_ (.I(_05321_),
    .Z(_05324_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10689_ (.I(_05309_),
    .Z(_05325_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10690_ (.A1(\soc.spi_video_ram_1.fifo_in_data[12] ),
    .A2(_05325_),
    .ZN(_05326_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10691_ (.A1(_03118_),
    .A2(_05324_),
    .B(_05326_),
    .ZN(_01258_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10692_ (.A1(\soc.spi_video_ram_1.fifo_in_data[13] ),
    .A2(_05325_),
    .ZN(_05327_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10693_ (.A1(_03202_),
    .A2(_05324_),
    .B(_05327_),
    .ZN(_01259_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10694_ (.A1(\soc.spi_video_ram_1.fifo_in_data[14] ),
    .A2(_05325_),
    .ZN(_05328_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10695_ (.A1(_03300_),
    .A2(_05324_),
    .B(_05328_),
    .ZN(_01260_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10696_ (.A1(\soc.spi_video_ram_1.fifo_in_data[15] ),
    .A2(_05325_),
    .ZN(_05329_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10697_ (.A1(_03396_),
    .A2(_05324_),
    .B(_05329_),
    .ZN(_01261_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10698_ (.I0(_02250_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[29][16] ),
    .S(_05321_),
    .Z(_05330_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10699_ (.I(_05330_),
    .Z(_01262_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10700_ (.I0(_02252_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[29][17] ),
    .S(_05321_),
    .Z(_05331_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10701_ (.I(_05331_),
    .Z(_01263_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10702_ (.I0(_02254_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[29][18] ),
    .S(_05321_),
    .Z(_05332_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10703_ (.I(_05332_),
    .Z(_01264_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10704_ (.I0(_02256_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[29][19] ),
    .S(_05321_),
    .Z(_05333_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10705_ (.I(_05333_),
    .Z(_01265_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10706_ (.I0(_02258_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[29][20] ),
    .S(_05321_),
    .Z(_05334_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10707_ (.I(_05334_),
    .Z(_01266_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10708_ (.A1(\soc.spi_video_ram_1.fifo_in_address[5] ),
    .A2(_05325_),
    .ZN(_05335_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10709_ (.A1(_03563_),
    .A2(_05324_),
    .B(_05335_),
    .ZN(_01267_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10710_ (.A1(\soc.spi_video_ram_1.fifo_in_address[6] ),
    .A2(_05325_),
    .ZN(_05336_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10711_ (.A1(_03494_),
    .A2(_05324_),
    .B(_05336_),
    .ZN(_01268_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10712_ (.A1(\soc.spi_video_ram_1.fifo_in_address[7] ),
    .A2(_05325_),
    .ZN(_05337_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10713_ (.A1(_03443_),
    .A2(_05324_),
    .B(_05337_),
    .ZN(_01269_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10714_ (.A1(\soc.spi_video_ram_1.fifo_in_address[8] ),
    .A2(_05325_),
    .ZN(_05338_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10715_ (.A1(_03347_),
    .A2(_05324_),
    .B(_05338_),
    .ZN(_01270_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10716_ (.A1(\soc.spi_video_ram_1.fifo_in_address[9] ),
    .A2(_05325_),
    .ZN(_05339_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10717_ (.A1(_03249_),
    .A2(_05324_),
    .B(_05339_),
    .ZN(_01271_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10718_ (.A1(\soc.spi_video_ram_1.fifo_in_address[10] ),
    .A2(_05325_),
    .ZN(_05340_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10719_ (.A1(_03160_),
    .A2(_05324_),
    .B(_05340_),
    .ZN(_01272_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10720_ (.I0(_02272_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[29][27] ),
    .S(_05321_),
    .Z(_05341_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10721_ (.I(_05341_),
    .Z(_01273_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10722_ (.I0(_02274_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[29][28] ),
    .S(_05321_),
    .Z(_05342_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10723_ (.I(_05342_),
    .Z(_01274_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10724_ (.A1(_01445_),
    .A2(_03931_),
    .Z(_05343_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _10725_ (.I(_05343_),
    .Z(_05344_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10726_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[31][0] ),
    .I1(\soc.spi_video_ram_1.fifo_in_data[0] ),
    .S(_05344_),
    .Z(_05345_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10727_ (.I(_05345_),
    .Z(_01275_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10728_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[31][1] ),
    .I1(\soc.spi_video_ram_1.fifo_in_data[1] ),
    .S(_05344_),
    .Z(_05346_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10729_ (.I(_05346_),
    .Z(_01276_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10730_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[31][2] ),
    .I1(\soc.spi_video_ram_1.fifo_in_data[2] ),
    .S(_05344_),
    .Z(_05347_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10731_ (.I(_05347_),
    .Z(_01277_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10732_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[31][3] ),
    .I1(\soc.spi_video_ram_1.fifo_in_data[3] ),
    .S(_05344_),
    .Z(_05348_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10733_ (.I(_05348_),
    .Z(_01278_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10734_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[31][4] ),
    .I1(\soc.spi_video_ram_1.fifo_in_data[4] ),
    .S(_05344_),
    .Z(_05349_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10735_ (.I(_05349_),
    .Z(_01279_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10736_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[31][5] ),
    .I1(\soc.spi_video_ram_1.fifo_in_data[5] ),
    .S(_05344_),
    .Z(_05350_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10737_ (.I(_05350_),
    .Z(_01280_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10738_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[31][6] ),
    .I1(\soc.spi_video_ram_1.fifo_in_data[6] ),
    .S(_05344_),
    .Z(_05351_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10739_ (.I(_05351_),
    .Z(_01281_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10740_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[31][7] ),
    .I1(\soc.spi_video_ram_1.fifo_in_data[7] ),
    .S(_05344_),
    .Z(_05352_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10741_ (.I(_05352_),
    .Z(_01282_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10742_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[31][8] ),
    .I1(\soc.spi_video_ram_1.fifo_in_data[8] ),
    .S(_05344_),
    .Z(_05353_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10743_ (.I(_05353_),
    .Z(_01283_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10744_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[31][9] ),
    .I1(\soc.spi_video_ram_1.fifo_in_data[9] ),
    .S(_05344_),
    .Z(_05354_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10745_ (.I(_05354_),
    .Z(_01284_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _10746_ (.I(_05343_),
    .Z(_05355_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10747_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[31][10] ),
    .I1(\soc.spi_video_ram_1.fifo_in_data[10] ),
    .S(_05355_),
    .Z(_05356_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10748_ (.I(_05356_),
    .Z(_01285_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10749_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[31][11] ),
    .I1(\soc.spi_video_ram_1.fifo_in_data[11] ),
    .S(_05355_),
    .Z(_05357_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10750_ (.I(_05357_),
    .Z(_01286_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10751_ (.I(_05355_),
    .Z(_05358_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10752_ (.I(_05343_),
    .Z(_05359_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10753_ (.A1(_04047_),
    .A2(_05359_),
    .ZN(_05360_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10754_ (.A1(_03121_),
    .A2(_05358_),
    .B(_05360_),
    .ZN(_01287_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10755_ (.A1(_04050_),
    .A2(_05359_),
    .ZN(_05361_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10756_ (.A1(_03199_),
    .A2(_05358_),
    .B(_05361_),
    .ZN(_01288_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10757_ (.A1(_04052_),
    .A2(_05359_),
    .ZN(_05362_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10758_ (.A1(_03297_),
    .A2(_05358_),
    .B(_05362_),
    .ZN(_01289_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10759_ (.A1(_04054_),
    .A2(_05359_),
    .ZN(_05363_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10760_ (.A1(_03393_),
    .A2(_05358_),
    .B(_05363_),
    .ZN(_01290_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10761_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[31][16] ),
    .I1(\soc.spi_video_ram_1.fifo_in_address[0] ),
    .S(_05355_),
    .Z(_05364_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10762_ (.I(_05364_),
    .Z(_01291_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10763_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[31][17] ),
    .I1(\soc.spi_video_ram_1.fifo_in_address[1] ),
    .S(_05355_),
    .Z(_05365_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10764_ (.I(_05365_),
    .Z(_01292_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10765_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[31][18] ),
    .I1(\soc.spi_video_ram_1.fifo_in_address[2] ),
    .S(_05355_),
    .Z(_05366_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10766_ (.I(_05366_),
    .Z(_01293_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10767_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[31][19] ),
    .I1(\soc.spi_video_ram_1.fifo_in_address[3] ),
    .S(_05355_),
    .Z(_05367_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10768_ (.I(_05367_),
    .Z(_01294_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10769_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[31][20] ),
    .I1(\soc.spi_video_ram_1.fifo_in_address[4] ),
    .S(_05355_),
    .Z(_05368_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10770_ (.I(_05368_),
    .Z(_01295_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10771_ (.A1(_04061_),
    .A2(_05359_),
    .ZN(_05369_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10772_ (.A1(_03566_),
    .A2(_05358_),
    .B(_05369_),
    .ZN(_01296_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10773_ (.A1(_04063_),
    .A2(_05359_),
    .ZN(_05370_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10774_ (.A1(_03491_),
    .A2(_05358_),
    .B(_05370_),
    .ZN(_01297_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10775_ (.A1(_04065_),
    .A2(_05359_),
    .ZN(_05371_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10776_ (.A1(_03440_),
    .A2(_05358_),
    .B(_05371_),
    .ZN(_01298_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10777_ (.A1(_04067_),
    .A2(_05359_),
    .ZN(_05372_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10778_ (.A1(_03344_),
    .A2(_05358_),
    .B(_05372_),
    .ZN(_01299_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10779_ (.A1(_04069_),
    .A2(_05359_),
    .ZN(_05373_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10780_ (.A1(_03246_),
    .A2(_05358_),
    .B(_05373_),
    .ZN(_01300_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10781_ (.A1(_03927_),
    .A2(_05359_),
    .ZN(_05374_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10782_ (.A1(_03157_),
    .A2(_05358_),
    .B(_05374_),
    .ZN(_01301_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10783_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[31][27] ),
    .I1(\soc.spi_video_ram_1.fifo_in_address[11] ),
    .S(_05355_),
    .Z(_05375_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10784_ (.I(_05375_),
    .Z(_01302_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10785_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[31][28] ),
    .I1(\soc.spi_video_ram_1.fifo_in_address[12] ),
    .S(_05355_),
    .Z(_05376_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10786_ (.I(_05376_),
    .Z(_01303_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _10787_ (.A1(_01445_),
    .A2(_04392_),
    .ZN(_05377_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _10788_ (.I(_05377_),
    .Z(_05378_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10789_ (.I0(_02213_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[7][0] ),
    .S(_05378_),
    .Z(_05379_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10790_ (.I(_05379_),
    .Z(_01304_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10791_ (.I0(_02219_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[7][1] ),
    .S(_05378_),
    .Z(_05380_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10792_ (.I(_05380_),
    .Z(_01305_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10793_ (.I0(_02221_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[7][2] ),
    .S(_05378_),
    .Z(_05381_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10794_ (.I(_05381_),
    .Z(_01306_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10795_ (.I0(_02223_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[7][3] ),
    .S(_05378_),
    .Z(_05382_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10796_ (.I(_05382_),
    .Z(_01307_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10797_ (.I0(_02225_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[7][4] ),
    .S(_05378_),
    .Z(_05383_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10798_ (.I(_05383_),
    .Z(_01308_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10799_ (.I0(_02227_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[7][5] ),
    .S(_05378_),
    .Z(_05384_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10800_ (.I(_05384_),
    .Z(_01309_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10801_ (.I0(_02229_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[7][6] ),
    .S(_05378_),
    .Z(_05385_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10802_ (.I(_05385_),
    .Z(_01310_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10803_ (.I0(_02231_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[7][7] ),
    .S(_05378_),
    .Z(_05386_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10804_ (.I(_05386_),
    .Z(_01311_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10805_ (.I0(_02233_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[7][8] ),
    .S(_05378_),
    .Z(_05387_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10806_ (.I(_05387_),
    .Z(_01312_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10807_ (.I0(_02235_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[7][9] ),
    .S(_05378_),
    .Z(_05388_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10808_ (.I(_05388_),
    .Z(_01313_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _10809_ (.I(_05377_),
    .Z(_05389_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10810_ (.I0(_02237_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[7][10] ),
    .S(_05389_),
    .Z(_05390_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10811_ (.I(_05390_),
    .Z(_01314_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10812_ (.I0(_02240_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[7][11] ),
    .S(_05389_),
    .Z(_05391_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10813_ (.I(_05391_),
    .Z(_01315_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10814_ (.I(_05389_),
    .Z(_05392_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10815_ (.I(_05377_),
    .Z(_05393_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10816_ (.A1(\soc.spi_video_ram_1.fifo_in_data[12] ),
    .A2(_05393_),
    .ZN(_05394_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10817_ (.A1(_03131_),
    .A2(_05392_),
    .B(_05394_),
    .ZN(_01316_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10818_ (.A1(\soc.spi_video_ram_1.fifo_in_data[13] ),
    .A2(_05393_),
    .ZN(_05395_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10819_ (.A1(_03222_),
    .A2(_05392_),
    .B(_05395_),
    .ZN(_01317_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10820_ (.A1(\soc.spi_video_ram_1.fifo_in_data[14] ),
    .A2(_05393_),
    .ZN(_05396_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10821_ (.A1(_03323_),
    .A2(_05392_),
    .B(_05396_),
    .ZN(_01318_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10822_ (.A1(\soc.spi_video_ram_1.fifo_in_data[15] ),
    .A2(_05393_),
    .ZN(_05397_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10823_ (.A1(_03416_),
    .A2(_05392_),
    .B(_05397_),
    .ZN(_01319_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10824_ (.I0(_02250_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[7][16] ),
    .S(_05389_),
    .Z(_05398_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10825_ (.I(_05398_),
    .Z(_01320_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10826_ (.I0(_02252_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[7][17] ),
    .S(_05389_),
    .Z(_05399_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10827_ (.I(_05399_),
    .Z(_01321_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10828_ (.I0(_02254_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[7][18] ),
    .S(_05389_),
    .Z(_05400_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10829_ (.I(_05400_),
    .Z(_01322_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10830_ (.I0(_02256_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[7][19] ),
    .S(_05389_),
    .Z(_05401_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10831_ (.I(_05401_),
    .Z(_01323_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10832_ (.I0(_02258_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[7][20] ),
    .S(_05389_),
    .Z(_05402_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10833_ (.I(_05402_),
    .Z(_01324_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10834_ (.A1(\soc.spi_video_ram_1.fifo_in_address[5] ),
    .A2(_05393_),
    .ZN(_05403_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10835_ (.A1(_03527_),
    .A2(_05392_),
    .B(_05403_),
    .ZN(_01325_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10836_ (.A1(\soc.spi_video_ram_1.fifo_in_address[6] ),
    .A2(_05393_),
    .ZN(_05404_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10837_ (.A1(_03501_),
    .A2(_05392_),
    .B(_05404_),
    .ZN(_01326_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10838_ (.A1(\soc.spi_video_ram_1.fifo_in_address[7] ),
    .A2(_05393_),
    .ZN(_05405_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10839_ (.A1(_03450_),
    .A2(_05392_),
    .B(_05405_),
    .ZN(_01327_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10840_ (.A1(\soc.spi_video_ram_1.fifo_in_address[8] ),
    .A2(_05393_),
    .ZN(_05406_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10841_ (.A1(_03354_),
    .A2(_05392_),
    .B(_05406_),
    .ZN(_01328_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10842_ (.A1(\soc.spi_video_ram_1.fifo_in_address[9] ),
    .A2(_05393_),
    .ZN(_05407_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10843_ (.A1(_03259_),
    .A2(_05392_),
    .B(_05407_),
    .ZN(_01329_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10844_ (.A1(\soc.spi_video_ram_1.fifo_in_address[10] ),
    .A2(_05393_),
    .ZN(_05408_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10845_ (.A1(_03175_),
    .A2(_05392_),
    .B(_05408_),
    .ZN(_01330_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10846_ (.I0(_02272_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[7][27] ),
    .S(_05389_),
    .Z(_05409_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10847_ (.I(_05409_),
    .Z(_01331_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10848_ (.I0(_02274_),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[7][28] ),
    .S(_05389_),
    .Z(_05410_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10849_ (.I(_05410_),
    .Z(_01332_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _10850_ (.A1(_05219_),
    .A2(_05244_),
    .ZN(_05411_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10851_ (.I(_05411_),
    .Z(_05412_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10852_ (.I(\soc.ram_encoder_0.data_out[0] ),
    .ZN(_05413_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _10853_ (.A1(_01589_),
    .A2(_05222_),
    .B1(_05412_),
    .B2(_05413_),
    .ZN(_01333_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10854_ (.I(\soc.ram_encoder_0.data_out[1] ),
    .ZN(_05414_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _10855_ (.A1(_01613_),
    .A2(_05222_),
    .B1(_05412_),
    .B2(_05414_),
    .ZN(_01334_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10856_ (.I(\soc.ram_encoder_0.data_out[2] ),
    .ZN(_05415_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _10857_ (.A1(_01632_),
    .A2(_05222_),
    .B1(_05412_),
    .B2(_05415_),
    .ZN(_01335_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10858_ (.I(\soc.ram_encoder_0.data_out[3] ),
    .ZN(_05416_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _10859_ (.A1(_01652_),
    .A2(_05222_),
    .B1(_05412_),
    .B2(_05416_),
    .ZN(_01336_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10860_ (.I(\soc.ram_encoder_0.data_out[4] ),
    .ZN(_05417_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _10861_ (.A1(_01666_),
    .A2(_05222_),
    .B1(_05412_),
    .B2(_05417_),
    .ZN(_01337_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10862_ (.I(\soc.ram_encoder_0.data_out[5] ),
    .ZN(_05418_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _10863_ (.A1(_01680_),
    .A2(_05222_),
    .B1(_05412_),
    .B2(_05418_),
    .ZN(_01338_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10864_ (.I(\soc.ram_encoder_0.data_out[6] ),
    .ZN(_05419_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _10865_ (.A1(_01699_),
    .A2(_05222_),
    .B1(_05412_),
    .B2(_05419_),
    .ZN(_01339_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10866_ (.I(\soc.ram_encoder_0.data_out[7] ),
    .ZN(_05420_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _10867_ (.A1(_01713_),
    .A2(_05222_),
    .B1(_05412_),
    .B2(_05420_),
    .ZN(_01340_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10868_ (.I(\soc.ram_encoder_0.data_out[8] ),
    .ZN(_05421_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _10869_ (.A1(_01736_),
    .A2(_05221_),
    .B1(_05412_),
    .B2(_05421_),
    .ZN(_01341_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10870_ (.I(\soc.ram_encoder_0.data_out[9] ),
    .ZN(_05422_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _10871_ (.A1(_01752_),
    .A2(_05221_),
    .B1(_05412_),
    .B2(_05422_),
    .ZN(_01342_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10872_ (.I(\soc.ram_encoder_0.data_out[10] ),
    .ZN(_05423_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _10873_ (.A1(_01767_),
    .A2(_05221_),
    .B1(_05411_),
    .B2(_05423_),
    .ZN(_01343_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10874_ (.I(\soc.ram_encoder_0.data_out[11] ),
    .ZN(_05424_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _10875_ (.A1(_01779_),
    .A2(_05221_),
    .B1(_05411_),
    .B2(_05424_),
    .ZN(_01344_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10876_ (.I(\soc.ram_encoder_0.data_out[12] ),
    .ZN(_05425_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _10877_ (.A1(_01803_),
    .A2(_05221_),
    .B1(_05411_),
    .B2(_05425_),
    .ZN(_01345_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10878_ (.I(\soc.ram_encoder_0.data_out[13] ),
    .ZN(_05426_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _10879_ (.A1(_01819_),
    .A2(_05221_),
    .B1(_05411_),
    .B2(_05426_),
    .ZN(_01346_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10880_ (.I(\soc.ram_encoder_0.data_out[14] ),
    .ZN(_05427_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _10881_ (.A1(_01834_),
    .A2(_05221_),
    .B1(_05411_),
    .B2(_05427_),
    .ZN(_01347_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10882_ (.I(\soc.ram_encoder_0.data_out[15] ),
    .ZN(_05428_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _10883_ (.A1(_02539_),
    .A2(_05221_),
    .B1(_05411_),
    .B2(_05428_),
    .ZN(_01348_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10884_ (.A1(_02214_),
    .A2(_03729_),
    .Z(_05429_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _10885_ (.I(_05429_),
    .Z(_05430_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _10886_ (.I(_05430_),
    .Z(_05431_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10887_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[8][0] ),
    .I1(\soc.spi_video_ram_1.fifo_in_data[0] ),
    .S(_05431_),
    .Z(_05432_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10888_ (.I(_05432_),
    .Z(_01349_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10889_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[8][1] ),
    .I1(\soc.spi_video_ram_1.fifo_in_data[1] ),
    .S(_05431_),
    .Z(_05433_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10890_ (.I(_05433_),
    .Z(_01350_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10891_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[8][2] ),
    .I1(\soc.spi_video_ram_1.fifo_in_data[2] ),
    .S(_05431_),
    .Z(_05434_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10892_ (.I(_05434_),
    .Z(_01351_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10893_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[8][3] ),
    .I1(\soc.spi_video_ram_1.fifo_in_data[3] ),
    .S(_05431_),
    .Z(_05435_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10894_ (.I(_05435_),
    .Z(_01352_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10895_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[8][4] ),
    .I1(\soc.spi_video_ram_1.fifo_in_data[4] ),
    .S(_05431_),
    .Z(_05436_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10896_ (.I(_05436_),
    .Z(_01353_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10897_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[8][5] ),
    .I1(\soc.spi_video_ram_1.fifo_in_data[5] ),
    .S(_05431_),
    .Z(_05437_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10898_ (.I(_05437_),
    .Z(_01354_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10899_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[8][6] ),
    .I1(\soc.spi_video_ram_1.fifo_in_data[6] ),
    .S(_05431_),
    .Z(_05438_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10900_ (.I(_05438_),
    .Z(_01355_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10901_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[8][7] ),
    .I1(\soc.spi_video_ram_1.fifo_in_data[7] ),
    .S(_05431_),
    .Z(_05439_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10902_ (.I(_05439_),
    .Z(_01356_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10903_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[8][8] ),
    .I1(\soc.spi_video_ram_1.fifo_in_data[8] ),
    .S(_05431_),
    .Z(_05440_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10904_ (.I(_05440_),
    .Z(_01357_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10905_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[8][9] ),
    .I1(\soc.spi_video_ram_1.fifo_in_data[9] ),
    .S(_05431_),
    .Z(_05441_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10906_ (.I(_05441_),
    .Z(_01358_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _10907_ (.I(_05429_),
    .Z(_05442_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10908_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[8][10] ),
    .I1(\soc.spi_video_ram_1.fifo_in_data[10] ),
    .S(_05442_),
    .Z(_05443_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10909_ (.I(_05443_),
    .Z(_01359_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10910_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[8][11] ),
    .I1(\soc.spi_video_ram_1.fifo_in_data[11] ),
    .S(_05442_),
    .Z(_05444_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10911_ (.I(_05444_),
    .Z(_01360_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10912_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[8][12] ),
    .I1(_04047_),
    .S(_05442_),
    .Z(_05445_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10913_ (.I(_05445_),
    .Z(_01361_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10914_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[8][13] ),
    .I1(_04050_),
    .S(_05442_),
    .Z(_05446_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10915_ (.I(_05446_),
    .Z(_01362_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10916_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[8][14] ),
    .I1(_04052_),
    .S(_05442_),
    .Z(_05447_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10917_ (.I(_05447_),
    .Z(_01363_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10918_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[8][15] ),
    .I1(_04054_),
    .S(_05442_),
    .Z(_05448_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10919_ (.I(_05448_),
    .Z(_01364_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10920_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[8][16] ),
    .I1(\soc.spi_video_ram_1.fifo_in_address[0] ),
    .S(_05442_),
    .Z(_05449_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10921_ (.I(_05449_),
    .Z(_01365_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10922_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[8][17] ),
    .I1(\soc.spi_video_ram_1.fifo_in_address[1] ),
    .S(_05442_),
    .Z(_05450_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10923_ (.I(_05450_),
    .Z(_01366_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10924_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[8][18] ),
    .I1(\soc.spi_video_ram_1.fifo_in_address[2] ),
    .S(_05442_),
    .Z(_05451_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10925_ (.I(_05451_),
    .Z(_01367_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10926_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[8][19] ),
    .I1(\soc.spi_video_ram_1.fifo_in_address[3] ),
    .S(_05442_),
    .Z(_05452_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10927_ (.I(_05452_),
    .Z(_01368_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10928_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[8][20] ),
    .I1(\soc.spi_video_ram_1.fifo_in_address[4] ),
    .S(_05430_),
    .Z(_05453_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10929_ (.I(_05453_),
    .Z(_01369_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10930_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[8][21] ),
    .I1(_04061_),
    .S(_05430_),
    .Z(_05454_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10931_ (.I(_05454_),
    .Z(_01370_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10932_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[8][22] ),
    .I1(_04063_),
    .S(_05430_),
    .Z(_05455_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10933_ (.I(_05455_),
    .Z(_01371_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10934_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[8][23] ),
    .I1(_04065_),
    .S(_05430_),
    .Z(_05456_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10935_ (.I(_05456_),
    .Z(_01372_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10936_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[8][24] ),
    .I1(_04067_),
    .S(_05430_),
    .Z(_05457_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10937_ (.I(_05457_),
    .Z(_01373_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10938_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[8][25] ),
    .I1(_04069_),
    .S(_05430_),
    .Z(_05458_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10939_ (.I(_05458_),
    .Z(_01374_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10940_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[8][26] ),
    .I1(_03927_),
    .S(_05430_),
    .Z(_05459_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10941_ (.I(_05459_),
    .Z(_01375_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10942_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[8][27] ),
    .I1(\soc.spi_video_ram_1.fifo_in_address[11] ),
    .S(_05430_),
    .Z(_05460_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10943_ (.I(_05460_),
    .Z(_01376_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10944_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[8][28] ),
    .I1(\soc.spi_video_ram_1.fifo_in_address[12] ),
    .S(_05430_),
    .Z(_05461_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10945_ (.I(_05461_),
    .Z(_01377_));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10946_ (.D(_00012_),
    .CLK(clknet_leaf_207_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[18][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10947_ (.D(_00013_),
    .CLK(clknet_leaf_216_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[18][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10948_ (.D(_00014_),
    .CLK(clknet_leaf_198_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[18][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10949_ (.D(_00015_),
    .CLK(clknet_leaf_140_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[18][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10950_ (.D(_00016_),
    .CLK(clknet_leaf_139_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[18][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10951_ (.D(_00017_),
    .CLK(clknet_leaf_215_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[18][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10952_ (.D(_00018_),
    .CLK(clknet_leaf_247_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[18][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10953_ (.D(_00019_),
    .CLK(clknet_leaf_194_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[18][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10954_ (.D(_00020_),
    .CLK(clknet_leaf_219_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[18][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10955_ (.D(_00021_),
    .CLK(clknet_leaf_255_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[18][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10956_ (.D(_00022_),
    .CLK(clknet_leaf_18_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[18][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10957_ (.D(_00023_),
    .CLK(clknet_leaf_33_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[18][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10958_ (.D(_00024_),
    .CLK(clknet_leaf_2_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[18][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10959_ (.D(_00025_),
    .CLK(clknet_leaf_40_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[18][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10960_ (.D(_00026_),
    .CLK(clknet_leaf_4_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[18][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10961_ (.D(_00027_),
    .CLK(clknet_leaf_10_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[18][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10962_ (.D(_00028_),
    .CLK(clknet_leaf_79_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[18][16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10963_ (.D(_00029_),
    .CLK(clknet_leaf_79_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[18][17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10964_ (.D(_00030_),
    .CLK(clknet_leaf_76_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[18][18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10965_ (.D(_00031_),
    .CLK(clknet_leaf_67_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[18][19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10966_ (.D(_00032_),
    .CLK(clknet_leaf_51_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[18][20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10967_ (.D(_00033_),
    .CLK(clknet_leaf_241_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[18][21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10968_ (.D(_00034_),
    .CLK(clknet_leaf_252_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[18][22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10969_ (.D(_00035_),
    .CLK(clknet_leaf_234_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[18][23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10970_ (.D(_00036_),
    .CLK(clknet_leaf_301_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[18][24] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10971_ (.D(_00037_),
    .CLK(clknet_leaf_234_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[18][25] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10972_ (.D(_00038_),
    .CLK(clknet_leaf_288_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[18][26] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10973_ (.D(_00039_),
    .CLK(clknet_leaf_271_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[18][27] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10974_ (.D(_00040_),
    .CLK(clknet_leaf_303_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[18][28] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10975_ (.D(_00041_),
    .CLK(clknet_5_23_0_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[17][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10976_ (.D(_00042_),
    .CLK(clknet_leaf_217_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[17][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10977_ (.D(_00043_),
    .CLK(clknet_leaf_197_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[17][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10978_ (.D(_00044_),
    .CLK(clknet_leaf_140_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[17][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10979_ (.D(_00045_),
    .CLK(clknet_leaf_140_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[17][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10980_ (.D(_00046_),
    .CLK(clknet_leaf_226_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[17][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10981_ (.D(_00047_),
    .CLK(clknet_leaf_211_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[17][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10982_ (.D(_00048_),
    .CLK(clknet_leaf_186_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[17][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10983_ (.D(_00049_),
    .CLK(clknet_5_23_0_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[17][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10984_ (.D(_00050_),
    .CLK(clknet_leaf_248_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[17][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10985_ (.D(_00051_),
    .CLK(clknet_leaf_13_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[17][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10986_ (.D(_00052_),
    .CLK(clknet_leaf_37_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[17][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10987_ (.D(_00053_),
    .CLK(clknet_leaf_2_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[17][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10988_ (.D(_00054_),
    .CLK(clknet_leaf_39_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[17][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10989_ (.D(_00055_),
    .CLK(clknet_leaf_4_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[17][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10990_ (.D(_00056_),
    .CLK(clknet_leaf_10_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[17][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10991_ (.D(_00057_),
    .CLK(clknet_leaf_76_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[17][16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10992_ (.D(_00058_),
    .CLK(clknet_leaf_79_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[17][17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10993_ (.D(_00059_),
    .CLK(clknet_leaf_76_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[17][18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10994_ (.D(_00060_),
    .CLK(clknet_leaf_68_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[17][19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10995_ (.D(_00061_),
    .CLK(clknet_leaf_264_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[17][20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10996_ (.D(_00062_),
    .CLK(clknet_leaf_235_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[17][21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10997_ (.D(_00063_),
    .CLK(clknet_leaf_267_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[17][22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10998_ (.D(_00064_),
    .CLK(clknet_leaf_233_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[17][23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _10999_ (.D(_00065_),
    .CLK(clknet_leaf_301_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[17][24] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11000_ (.D(_00066_),
    .CLK(clknet_leaf_235_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[17][25] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11001_ (.D(_00067_),
    .CLK(clknet_leaf_288_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[17][26] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11002_ (.D(_00068_),
    .CLK(clknet_leaf_265_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[17][27] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11003_ (.D(_00069_),
    .CLK(clknet_leaf_278_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[17][28] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11004_ (.D(_00070_),
    .CLK(clknet_leaf_222_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[16][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11005_ (.D(_00071_),
    .CLK(clknet_leaf_218_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[16][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11006_ (.D(_00072_),
    .CLK(clknet_leaf_197_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[16][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11007_ (.D(_00073_),
    .CLK(clknet_leaf_138_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[16][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11008_ (.D(_00074_),
    .CLK(clknet_leaf_140_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[16][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11009_ (.D(_00075_),
    .CLK(clknet_leaf_217_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[16][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11010_ (.D(_00076_),
    .CLK(clknet_leaf_211_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[16][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11011_ (.D(_00077_),
    .CLK(clknet_leaf_187_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[16][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11012_ (.D(_00078_),
    .CLK(clknet_leaf_218_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[16][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11013_ (.D(_00079_),
    .CLK(clknet_leaf_248_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[16][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11014_ (.D(_00080_),
    .CLK(clknet_leaf_13_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[16][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11015_ (.D(_00081_),
    .CLK(clknet_leaf_42_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[16][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11016_ (.D(_00082_),
    .CLK(clknet_leaf_4_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[16][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11017_ (.D(_00083_),
    .CLK(clknet_leaf_11_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[16][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11018_ (.D(_00084_),
    .CLK(clknet_leaf_4_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[16][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11019_ (.D(_00085_),
    .CLK(clknet_leaf_10_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[16][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11020_ (.D(_00086_),
    .CLK(clknet_leaf_75_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[16][16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11021_ (.D(_00087_),
    .CLK(clknet_leaf_80_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[16][17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11022_ (.D(_00088_),
    .CLK(clknet_leaf_75_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[16][18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11023_ (.D(_00089_),
    .CLK(clknet_leaf_67_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[16][19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11024_ (.D(_00090_),
    .CLK(clknet_leaf_263_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[16][20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11025_ (.D(_00091_),
    .CLK(clknet_leaf_236_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[16][21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11026_ (.D(_00092_),
    .CLK(clknet_leaf_266_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[16][22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11027_ (.D(_00093_),
    .CLK(clknet_leaf_236_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[16][23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11028_ (.D(_00094_),
    .CLK(clknet_leaf_304_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[16][24] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11029_ (.D(_00095_),
    .CLK(clknet_leaf_236_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[16][25] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11030_ (.D(_00096_),
    .CLK(clknet_leaf_287_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[16][26] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11031_ (.D(_00097_),
    .CLK(clknet_leaf_271_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[16][27] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11032_ (.D(_00098_),
    .CLK(clknet_leaf_277_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[16][28] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11033_ (.D(_00099_),
    .CLK(clknet_leaf_219_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[0][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11034_ (.D(_00100_),
    .CLK(clknet_leaf_215_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[0][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11035_ (.D(_00101_),
    .CLK(clknet_leaf_257_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[0][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11036_ (.D(_00102_),
    .CLK(clknet_leaf_199_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[0][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11037_ (.D(_00103_),
    .CLK(clknet_leaf_200_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[0][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11038_ (.D(_00104_),
    .CLK(clknet_leaf_226_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[0][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11039_ (.D(_00105_),
    .CLK(clknet_leaf_247_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[0][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11040_ (.D(_00106_),
    .CLK(clknet_leaf_205_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[0][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11041_ (.D(_00107_),
    .CLK(clknet_leaf_220_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[0][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11042_ (.D(_00108_),
    .CLK(clknet_leaf_247_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[0][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11043_ (.D(_00109_),
    .CLK(clknet_leaf_18_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[0][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11044_ (.D(_00110_),
    .CLK(clknet_leaf_36_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[0][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11045_ (.D(_00111_),
    .CLK(clknet_leaf_0_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[0][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11046_ (.D(_00112_),
    .CLK(clknet_leaf_320_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[0][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11047_ (.D(_00113_),
    .CLK(clknet_leaf_321_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[0][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11048_ (.D(_00114_),
    .CLK(clknet_leaf_321_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[0][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11049_ (.D(_00115_),
    .CLK(clknet_leaf_77_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[0][16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11050_ (.D(_00116_),
    .CLK(clknet_leaf_78_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[0][17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11051_ (.D(_00117_),
    .CLK(clknet_leaf_76_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[0][18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11052_ (.D(_00118_),
    .CLK(clknet_leaf_70_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[0][19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11053_ (.D(_00119_),
    .CLK(clknet_leaf_51_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[0][20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11054_ (.D(_00120_),
    .CLK(clknet_leaf_229_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[0][21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11055_ (.D(_00121_),
    .CLK(clknet_leaf_249_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[0][22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11056_ (.D(_00122_),
    .CLK(clknet_leaf_242_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[0][23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11057_ (.D(_00123_),
    .CLK(clknet_leaf_296_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[0][24] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11058_ (.D(_00124_),
    .CLK(clknet_leaf_229_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[0][25] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11059_ (.D(_00125_),
    .CLK(clknet_leaf_293_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[0][26] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11060_ (.D(_00126_),
    .CLK(clknet_leaf_43_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[0][27] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11061_ (.D(_00127_),
    .CLK(clknet_leaf_296_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[0][28] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11062_ (.D(_00128_),
    .CLK(clknet_leaf_177_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[13][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11063_ (.D(_00129_),
    .CLK(clknet_leaf_224_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[13][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11064_ (.D(_00130_),
    .CLK(clknet_leaf_137_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[13][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11065_ (.D(_00131_),
    .CLK(clknet_leaf_262_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[13][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11066_ (.D(_00132_),
    .CLK(clknet_leaf_260_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[13][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11067_ (.D(_00133_),
    .CLK(clknet_leaf_219_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[13][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11068_ (.D(_00134_),
    .CLK(clknet_leaf_208_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[13][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11069_ (.D(_00135_),
    .CLK(clknet_leaf_191_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[13][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11070_ (.D(_00136_),
    .CLK(clknet_leaf_176_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[13][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11071_ (.D(_00137_),
    .CLK(clknet_leaf_202_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[13][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11072_ (.D(_00138_),
    .CLK(clknet_leaf_16_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[13][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11073_ (.D(_00139_),
    .CLK(clknet_leaf_38_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[13][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11074_ (.D(_00140_),
    .CLK(clknet_leaf_7_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[13][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11075_ (.D(_00141_),
    .CLK(clknet_leaf_16_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[13][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11076_ (.D(_00142_),
    .CLK(clknet_leaf_5_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[13][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11077_ (.D(_00143_),
    .CLK(clknet_leaf_3_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[13][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11078_ (.D(_00144_),
    .CLK(clknet_leaf_20_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[13][16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11079_ (.D(_00145_),
    .CLK(clknet_leaf_20_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[13][17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11080_ (.D(_00146_),
    .CLK(clknet_leaf_21_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[13][18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11081_ (.D(_00147_),
    .CLK(clknet_leaf_35_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[13][19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11082_ (.D(_00148_),
    .CLK(clknet_leaf_48_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[13][20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11083_ (.D(_00149_),
    .CLK(clknet_leaf_283_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[13][21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11084_ (.D(_00150_),
    .CLK(clknet_leaf_267_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[13][22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11085_ (.D(_00151_),
    .CLK(clknet_leaf_285_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[13][23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11086_ (.D(_00152_),
    .CLK(clknet_leaf_305_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[13][24] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11087_ (.D(_00153_),
    .CLK(clknet_leaf_285_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[13][25] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11088_ (.D(_00154_),
    .CLK(clknet_leaf_279_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[13][26] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11089_ (.D(_00155_),
    .CLK(clknet_leaf_41_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[13][27] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11090_ (.D(_00156_),
    .CLK(clknet_leaf_282_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[13][28] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11091_ (.D(_00157_),
    .CLK(clknet_leaf_177_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[12][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11092_ (.D(_00158_),
    .CLK(clknet_leaf_224_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[12][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11093_ (.D(_00159_),
    .CLK(clknet_leaf_54_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[12][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11094_ (.D(_00160_),
    .CLK(clknet_leaf_261_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[12][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11095_ (.D(_00161_),
    .CLK(clknet_leaf_260_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[12][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11096_ (.D(_00162_),
    .CLK(clknet_leaf_224_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[12][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11097_ (.D(_00163_),
    .CLK(clknet_leaf_203_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[12][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11098_ (.D(_00164_),
    .CLK(clknet_leaf_205_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[12][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11099_ (.D(_00165_),
    .CLK(clknet_leaf_175_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[12][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11100_ (.D(_00166_),
    .CLK(clknet_leaf_202_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[12][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11101_ (.D(_00167_),
    .CLK(clknet_leaf_16_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[12][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11102_ (.D(_00168_),
    .CLK(clknet_leaf_38_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[12][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11103_ (.D(_00169_),
    .CLK(clknet_leaf_7_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[12][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11104_ (.D(_00170_),
    .CLK(clknet_leaf_16_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[12][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11105_ (.D(_00171_),
    .CLK(clknet_leaf_5_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[12][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11106_ (.D(_00172_),
    .CLK(clknet_leaf_3_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[12][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11107_ (.D(_00173_),
    .CLK(clknet_leaf_21_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[12][16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11108_ (.D(_00174_),
    .CLK(clknet_leaf_21_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[12][17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11109_ (.D(_00175_),
    .CLK(clknet_leaf_28_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[12][18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11110_ (.D(_00176_),
    .CLK(clknet_leaf_31_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[12][19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11111_ (.D(_00177_),
    .CLK(clknet_leaf_50_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[12][20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11112_ (.D(_00178_),
    .CLK(clknet_leaf_285_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[12][21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11113_ (.D(_00179_),
    .CLK(clknet_leaf_267_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[12][22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11114_ (.D(_00180_),
    .CLK(clknet_leaf_236_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[12][23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11115_ (.D(_00181_),
    .CLK(clknet_leaf_304_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[12][24] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11116_ (.D(_00182_),
    .CLK(clknet_leaf_286_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[12][25] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11117_ (.D(_00183_),
    .CLK(clknet_leaf_279_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[12][26] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11118_ (.D(_00184_),
    .CLK(clknet_leaf_43_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[12][27] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11119_ (.D(_00185_),
    .CLK(clknet_leaf_281_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[12][28] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11120_ (.D(_00186_),
    .CLK(clknet_leaf_178_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[14][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11121_ (.D(_00187_),
    .CLK(clknet_leaf_222_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[14][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11122_ (.D(_00188_),
    .CLK(clknet_leaf_54_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[14][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11123_ (.D(_00189_),
    .CLK(clknet_leaf_54_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[14][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11124_ (.D(_00190_),
    .CLK(clknet_leaf_54_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[14][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11125_ (.D(_00191_),
    .CLK(clknet_leaf_221_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[14][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11126_ (.D(_00192_),
    .CLK(clknet_leaf_202_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[14][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11127_ (.D(_00193_),
    .CLK(clknet_leaf_192_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[14][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11128_ (.D(_00194_),
    .CLK(clknet_leaf_176_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[14][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11129_ (.D(_00195_),
    .CLK(clknet_leaf_201_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[14][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11130_ (.D(_00196_),
    .CLK(clknet_leaf_16_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[14][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11131_ (.D(_00197_),
    .CLK(clknet_leaf_46_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[14][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11132_ (.D(_00198_),
    .CLK(clknet_leaf_310_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[14][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11133_ (.D(_00199_),
    .CLK(clknet_leaf_11_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[14][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11134_ (.D(_00200_),
    .CLK(clknet_leaf_310_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[14][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11135_ (.D(_00201_),
    .CLK(clknet_leaf_8_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[14][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11136_ (.D(_00202_),
    .CLK(clknet_leaf_20_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[14][16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11137_ (.D(_00203_),
    .CLK(clknet_leaf_22_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[14][17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11138_ (.D(_00204_),
    .CLK(clknet_leaf_22_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[14][18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11139_ (.D(_00205_),
    .CLK(clknet_leaf_28_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[14][19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11140_ (.D(_00206_),
    .CLK(clknet_leaf_48_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[14][20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11141_ (.D(_00207_),
    .CLK(clknet_leaf_282_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[14][21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11142_ (.D(_00208_),
    .CLK(clknet_leaf_268_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[14][22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11143_ (.D(_00209_),
    .CLK(clknet_leaf_284_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[14][23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11144_ (.D(_00210_),
    .CLK(clknet_leaf_306_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[14][24] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11145_ (.D(_00211_),
    .CLK(clknet_leaf_285_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[14][25] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11146_ (.D(_00212_),
    .CLK(clknet_leaf_278_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[14][26] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11147_ (.D(_00213_),
    .CLK(clknet_leaf_45_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[14][27] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11148_ (.D(_00214_),
    .CLK(clknet_leaf_282_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[14][28] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11149_ (.D(_00215_),
    .CLK(clknet_leaf_125_wb_clk_i),
    .Q(net65));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11150_ (.D(_00216_),
    .CLK(clknet_leaf_125_wb_clk_i),
    .Q(net66));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11151_ (.D(_00217_),
    .CLK(clknet_leaf_126_wb_clk_i),
    .Q(net67));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11152_ (.D(_00218_),
    .CLK(clknet_leaf_166_wb_clk_i),
    .Q(\soc.ram_encoder_0.output_bits_left[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11153_ (.D(_00219_),
    .CLK(clknet_leaf_166_wb_clk_i),
    .Q(\soc.ram_encoder_0.output_bits_left[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11154_ (.D(_00220_),
    .CLK(clknet_leaf_165_wb_clk_i),
    .Q(\soc.ram_encoder_0.output_bits_left[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11155_ (.D(_00221_),
    .CLK(clknet_leaf_95_wb_clk_i),
    .Q(\soc.rom_encoder_0.output_bits_left[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11156_ (.D(_00222_),
    .CLK(clknet_leaf_93_wb_clk_i),
    .Q(\soc.rom_encoder_0.output_bits_left[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11157_ (.D(_00223_),
    .CLK(clknet_leaf_95_wb_clk_i),
    .Q(\soc.rom_encoder_0.output_bits_left[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11158_ (.D(_00224_),
    .CLK(net84),
    .Q(\soc.cpu.AReg.data[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11159_ (.D(_00225_),
    .CLK(clknet_leaf_105_wb_clk_i),
    .Q(\soc.rom_encoder_0.output_buffer[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11160_ (.D(_00226_),
    .CLK(clknet_leaf_92_wb_clk_i),
    .Q(\soc.rom_encoder_0.output_buffer[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11161_ (.D(_00227_),
    .CLK(clknet_leaf_105_wb_clk_i),
    .Q(\soc.rom_encoder_0.output_buffer[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11162_ (.D(_00228_),
    .CLK(clknet_leaf_92_wb_clk_i),
    .Q(\soc.rom_encoder_0.output_buffer[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11163_ (.D(_00229_),
    .CLK(clknet_leaf_149_wb_clk_i),
    .Q(\soc.ram_encoder_0.output_buffer[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11164_ (.D(_00230_),
    .CLK(clknet_leaf_149_wb_clk_i),
    .Q(\soc.ram_encoder_0.output_buffer[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11165_ (.D(_00231_),
    .CLK(clknet_leaf_149_wb_clk_i),
    .Q(\soc.ram_encoder_0.output_buffer[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11166_ (.D(_00232_),
    .CLK(clknet_leaf_149_wb_clk_i),
    .Q(\soc.ram_encoder_0.output_buffer[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11167_ (.D(_00233_),
    .CLK(clknet_leaf_56_wb_clk_i),
    .Q(\soc.spi_video_ram_1.output_buffer[23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11168_ (.D(_00234_),
    .CLK(clknet_leaf_56_wb_clk_i),
    .Q(\soc.spi_video_ram_1.output_buffer[22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11169_ (.D(_00235_),
    .CLK(clknet_leaf_55_wb_clk_i),
    .Q(\soc.spi_video_ram_1.output_buffer[21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11170_ (.D(_00236_),
    .CLK(clknet_leaf_136_wb_clk_i),
    .Q(\soc.spi_video_ram_1.output_buffer[20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11171_ (.D(_00237_),
    .CLK(clknet_leaf_134_wb_clk_i),
    .Q(\soc.spi_video_ram_1.output_buffer[19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11172_ (.D(_00238_),
    .CLK(clknet_leaf_55_wb_clk_i),
    .Q(\soc.spi_video_ram_1.output_buffer[18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11173_ (.D(_00239_),
    .CLK(clknet_leaf_56_wb_clk_i),
    .Q(\soc.spi_video_ram_1.output_buffer[17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11174_ (.D(_00240_),
    .CLK(clknet_5_24_0_wb_clk_i),
    .Q(\soc.spi_video_ram_1.output_buffer[16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11175_ (.D(_00241_),
    .CLK(clknet_leaf_56_wb_clk_i),
    .Q(\soc.spi_video_ram_1.output_buffer[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11176_ (.D(_00242_),
    .CLK(clknet_leaf_56_wb_clk_i),
    .Q(\soc.spi_video_ram_1.output_buffer[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11177_ (.D(_00243_),
    .CLK(clknet_leaf_60_wb_clk_i),
    .Q(\soc.spi_video_ram_1.output_buffer[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11178_ (.D(_00244_),
    .CLK(clknet_leaf_60_wb_clk_i),
    .Q(\soc.spi_video_ram_1.output_buffer[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11179_ (.D(_00245_),
    .CLK(clknet_leaf_60_wb_clk_i),
    .Q(\soc.spi_video_ram_1.output_buffer[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11180_ (.D(_00246_),
    .CLK(clknet_leaf_58_wb_clk_i),
    .Q(\soc.spi_video_ram_1.output_buffer[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11181_ (.D(_00247_),
    .CLK(clknet_leaf_62_wb_clk_i),
    .Q(\soc.spi_video_ram_1.output_buffer[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11182_ (.D(_00248_),
    .CLK(clknet_leaf_62_wb_clk_i),
    .Q(\soc.spi_video_ram_1.output_buffer[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11183_ (.D(_00249_),
    .CLK(clknet_leaf_59_wb_clk_i),
    .Q(\soc.spi_video_ram_1.output_buffer[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11184_ (.D(_00250_),
    .CLK(clknet_leaf_56_wb_clk_i),
    .Q(\soc.spi_video_ram_1.output_buffer[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11185_ (.D(_00251_),
    .CLK(clknet_leaf_59_wb_clk_i),
    .Q(\soc.spi_video_ram_1.output_buffer[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11186_ (.D(_00252_),
    .CLK(clknet_leaf_58_wb_clk_i),
    .Q(\soc.spi_video_ram_1.output_buffer[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11187_ (.D(_00253_),
    .CLK(clknet_leaf_58_wb_clk_i),
    .Q(\soc.spi_video_ram_1.output_buffer[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11188_ (.D(_00254_),
    .CLK(clknet_leaf_60_wb_clk_i),
    .Q(\soc.spi_video_ram_1.output_buffer[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11189_ (.D(_00255_),
    .CLK(clknet_leaf_60_wb_clk_i),
    .Q(\soc.spi_video_ram_1.output_buffer[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11190_ (.D(_00256_),
    .CLK(clknet_leaf_191_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[11][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11191_ (.D(_00257_),
    .CLK(clknet_leaf_190_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[11][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11192_ (.D(_00258_),
    .CLK(clknet_leaf_137_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[11][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11193_ (.D(_00259_),
    .CLK(clknet_leaf_260_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[11][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11194_ (.D(_00260_),
    .CLK(clknet_leaf_196_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[11][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11195_ (.D(_00261_),
    .CLK(clknet_leaf_207_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[11][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11196_ (.D(_00262_),
    .CLK(clknet_leaf_203_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[11][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11197_ (.D(_00263_),
    .CLK(clknet_leaf_192_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[11][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11198_ (.D(_00264_),
    .CLK(clknet_leaf_189_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[11][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11199_ (.D(_00265_),
    .CLK(clknet_leaf_256_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[11][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11200_ (.D(_00266_),
    .CLK(clknet_leaf_15_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[11][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11201_ (.D(_00267_),
    .CLK(clknet_leaf_46_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[11][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11202_ (.D(_00268_),
    .CLK(clknet_leaf_2_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[11][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11203_ (.D(_00269_),
    .CLK(clknet_leaf_12_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[11][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11204_ (.D(_00270_),
    .CLK(clknet_leaf_5_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[11][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11205_ (.D(_00271_),
    .CLK(clknet_leaf_8_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[11][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11206_ (.D(_00272_),
    .CLK(clknet_leaf_26_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[11][16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11207_ (.D(_00273_),
    .CLK(clknet_leaf_24_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[11][17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11208_ (.D(_00274_),
    .CLK(clknet_leaf_25_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[11][18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11209_ (.D(_00275_),
    .CLK(clknet_leaf_30_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[11][19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11210_ (.D(_00276_),
    .CLK(clknet_leaf_52_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[11][20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11211_ (.D(_00277_),
    .CLK(clknet_leaf_282_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[11][21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11212_ (.D(_00278_),
    .CLK(clknet_leaf_254_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[11][22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11213_ (.D(_00279_),
    .CLK(clknet_leaf_238_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[11][23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11214_ (.D(_00280_),
    .CLK(clknet_leaf_304_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[11][24] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11215_ (.D(_00281_),
    .CLK(clknet_leaf_236_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[11][25] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11216_ (.D(_00282_),
    .CLK(clknet_leaf_280_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[11][26] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11217_ (.D(_00283_),
    .CLK(clknet_leaf_264_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[11][27] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11218_ (.D(_00284_),
    .CLK(clknet_leaf_269_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[11][28] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11219_ (.D(_00285_),
    .CLK(clknet_leaf_81_wb_clk_i),
    .Q(\soc.display_clks_before_active[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11220_ (.D(_00286_),
    .CLK(clknet_5_10_0_wb_clk_i),
    .Q(\soc.video_generator_1.h_count[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11221_ (.D(_00287_),
    .CLK(clknet_leaf_81_wb_clk_i),
    .Q(\soc.video_generator_1.h_count[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11222_ (.D(_00288_),
    .CLK(clknet_leaf_87_wb_clk_i),
    .Q(\soc.video_generator_1.h_count[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11223_ (.D(_00289_),
    .CLK(clknet_leaf_87_wb_clk_i),
    .Q(\soc.video_generator_1.h_count[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11224_ (.D(_00290_),
    .CLK(clknet_leaf_86_wb_clk_i),
    .Q(\soc.video_generator_1.h_count[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11225_ (.D(_00291_),
    .CLK(clknet_leaf_87_wb_clk_i),
    .Q(\soc.video_generator_1.h_count[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11226_ (.D(_00292_),
    .CLK(clknet_leaf_86_wb_clk_i),
    .Q(\soc.video_generator_1.h_count[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11227_ (.D(_00293_),
    .CLK(clknet_leaf_85_wb_clk_i),
    .Q(\soc.video_generator_1.h_count[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11228_ (.D(_00294_),
    .CLK(clknet_leaf_86_wb_clk_i),
    .Q(\soc.video_generator_1.h_count[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11229_ (.D(_00295_),
    .CLK(clknet_leaf_191_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[10][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11230_ (.D(_00296_),
    .CLK(clknet_leaf_205_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[10][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11231_ (.D(_00297_),
    .CLK(clknet_leaf_137_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[10][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11232_ (.D(_00298_),
    .CLK(clknet_leaf_260_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[10][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11233_ (.D(_00299_),
    .CLK(clknet_leaf_198_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[10][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11234_ (.D(_00300_),
    .CLK(clknet_leaf_205_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[10][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11235_ (.D(_00301_),
    .CLK(clknet_leaf_203_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[10][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11236_ (.D(_00302_),
    .CLK(clknet_leaf_192_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[10][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11237_ (.D(_00303_),
    .CLK(clknet_leaf_190_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[10][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11238_ (.D(_00304_),
    .CLK(clknet_leaf_256_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[10][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11239_ (.D(_00305_),
    .CLK(clknet_leaf_13_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[10][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11240_ (.D(_00306_),
    .CLK(clknet_leaf_38_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[10][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11241_ (.D(_00307_),
    .CLK(clknet_leaf_1_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[10][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11242_ (.D(_00308_),
    .CLK(clknet_leaf_12_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[10][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11243_ (.D(_00309_),
    .CLK(clknet_leaf_6_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[10][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11244_ (.D(_00310_),
    .CLK(clknet_leaf_3_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[10][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11245_ (.D(_00311_),
    .CLK(clknet_leaf_25_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[10][16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11246_ (.D(_00312_),
    .CLK(clknet_leaf_24_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[10][17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11247_ (.D(_00313_),
    .CLK(clknet_leaf_25_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[10][18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11248_ (.D(_00314_),
    .CLK(clknet_leaf_30_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[10][19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11249_ (.D(_00315_),
    .CLK(clknet_leaf_52_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[10][20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11250_ (.D(_00316_),
    .CLK(clknet_leaf_285_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[10][21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11251_ (.D(_00317_),
    .CLK(clknet_leaf_252_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[10][22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11252_ (.D(_00318_),
    .CLK(clknet_leaf_237_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[10][23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11253_ (.D(_00319_),
    .CLK(clknet_leaf_304_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[10][24] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11254_ (.D(_00320_),
    .CLK(clknet_leaf_236_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[10][25] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11255_ (.D(_00321_),
    .CLK(clknet_leaf_280_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[10][26] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11256_ (.D(_00322_),
    .CLK(clknet_leaf_271_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[10][27] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11257_ (.D(_00323_),
    .CLK(clknet_leaf_282_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[10][28] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11258_ (.D(_00324_),
    .CLK(clknet_leaf_99_wb_clk_i),
    .Q(net64));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11259_ (.D(_00325_),
    .CLK(clknet_leaf_149_wb_clk_i),
    .Q(\soc.ram_encoder_0.output_buffer[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11260_ (.D(_00326_),
    .CLK(clknet_leaf_150_wb_clk_i),
    .Q(\soc.ram_encoder_0.output_buffer[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11261_ (.D(_00327_),
    .CLK(clknet_leaf_150_wb_clk_i),
    .Q(\soc.ram_encoder_0.output_buffer[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11262_ (.D(_00328_),
    .CLK(clknet_leaf_151_wb_clk_i),
    .Q(\soc.ram_encoder_0.output_buffer[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11263_ (.D(_00329_),
    .CLK(clknet_leaf_151_wb_clk_i),
    .Q(\soc.ram_encoder_0.output_buffer[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11264_ (.D(_00330_),
    .CLK(clknet_leaf_169_wb_clk_i),
    .Q(\soc.ram_encoder_0.output_buffer[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11265_ (.D(_00331_),
    .CLK(clknet_leaf_169_wb_clk_i),
    .Q(\soc.ram_encoder_0.output_buffer[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11266_ (.D(_00332_),
    .CLK(clknet_leaf_168_wb_clk_i),
    .Q(\soc.ram_encoder_0.output_buffer[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11267_ (.D(_00333_),
    .CLK(clknet_leaf_168_wb_clk_i),
    .Q(\soc.ram_encoder_0.output_buffer[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11268_ (.D(_00334_),
    .CLK(clknet_leaf_167_wb_clk_i),
    .Q(\soc.ram_encoder_0.output_buffer[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11269_ (.D(_00335_),
    .CLK(clknet_leaf_167_wb_clk_i),
    .Q(\soc.ram_encoder_0.output_buffer[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11270_ (.D(_00336_),
    .CLK(clknet_leaf_167_wb_clk_i),
    .Q(\soc.ram_encoder_0.output_buffer[16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11271_ (.D(_00337_),
    .CLK(clknet_leaf_166_wb_clk_i),
    .Q(\soc.ram_encoder_0.output_buffer[17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11272_ (.D(_00338_),
    .CLK(clknet_leaf_166_wb_clk_i),
    .Q(\soc.ram_encoder_0.output_buffer[18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11273_ (.D(_00339_),
    .CLK(clknet_leaf_168_wb_clk_i),
    .Q(\soc.ram_encoder_0.output_buffer[19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11274_ (.D(_00340_),
    .CLK(clknet_leaf_221_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[1][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11275_ (.D(_00341_),
    .CLK(clknet_leaf_216_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[1][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11276_ (.D(_00342_),
    .CLK(clknet_leaf_258_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[1][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11277_ (.D(_00343_),
    .CLK(clknet_leaf_259_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[1][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11278_ (.D(_00344_),
    .CLK(clknet_leaf_200_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[1][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11279_ (.D(_00345_),
    .CLK(clknet_leaf_215_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[1][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11280_ (.D(_00346_),
    .CLK(clknet_leaf_213_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[1][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11281_ (.D(_00347_),
    .CLK(clknet_leaf_205_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[1][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11282_ (.D(_00348_),
    .CLK(clknet_leaf_220_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[1][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11283_ (.D(_00349_),
    .CLK(clknet_leaf_248_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[1][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11284_ (.D(_00350_),
    .CLK(clknet_leaf_17_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[1][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11285_ (.D(_00351_),
    .CLK(clknet_leaf_14_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[1][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11286_ (.D(_00352_),
    .CLK(clknet_leaf_0_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[1][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11287_ (.D(_00353_),
    .CLK(clknet_leaf_319_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[1][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11288_ (.D(_00354_),
    .CLK(clknet_leaf_317_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[1][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11289_ (.D(_00355_),
    .CLK(clknet_leaf_0_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[1][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11290_ (.D(_00356_),
    .CLK(clknet_leaf_77_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[1][16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11291_ (.D(_00357_),
    .CLK(clknet_leaf_78_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[1][17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11292_ (.D(_00358_),
    .CLK(clknet_leaf_77_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[1][18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11293_ (.D(_00359_),
    .CLK(clknet_leaf_68_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[1][19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11294_ (.D(_00360_),
    .CLK(clknet_leaf_44_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[1][20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11295_ (.D(_00361_),
    .CLK(clknet_leaf_229_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[1][21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11296_ (.D(_00362_),
    .CLK(clknet_leaf_251_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[1][22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11297_ (.D(_00363_),
    .CLK(clknet_leaf_242_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[1][23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11298_ (.D(_00364_),
    .CLK(clknet_leaf_296_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[1][24] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11299_ (.D(_00365_),
    .CLK(clknet_leaf_229_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[1][25] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11300_ (.D(_00366_),
    .CLK(clknet_leaf_293_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[1][26] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11301_ (.D(_00367_),
    .CLK(clknet_leaf_43_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[1][27] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11302_ (.D(_00368_),
    .CLK(clknet_leaf_297_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[1][28] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11303_ (.D(_00369_),
    .CLK(clknet_leaf_184_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[26][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11304_ (.D(_00370_),
    .CLK(clknet_leaf_187_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[26][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11305_ (.D(_00371_),
    .CLK(clknet_leaf_196_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[26][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11306_ (.D(_00372_),
    .CLK(clknet_leaf_142_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[26][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11307_ (.D(_00373_),
    .CLK(clknet_leaf_141_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[26][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11308_ (.D(_00374_),
    .CLK(clknet_leaf_188_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[26][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11309_ (.D(_00375_),
    .CLK(clknet_leaf_201_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[26][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11310_ (.D(_00376_),
    .CLK(clknet_leaf_146_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[26][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11311_ (.D(_00377_),
    .CLK(clknet_leaf_184_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[26][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11312_ (.D(_00378_),
    .CLK(clknet_leaf_259_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[26][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11313_ (.D(_00379_),
    .CLK(clknet_leaf_17_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[26][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11314_ (.D(_00380_),
    .CLK(clknet_leaf_34_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[26][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11315_ (.D(_00381_),
    .CLK(clknet_leaf_1_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[26][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11316_ (.D(_00382_),
    .CLK(clknet_leaf_315_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[26][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11317_ (.D(_00383_),
    .CLK(clknet_leaf_318_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[26][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11318_ (.D(_00384_),
    .CLK(clknet_leaf_314_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[26][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11319_ (.D(_00385_),
    .CLK(clknet_leaf_19_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[26][16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11320_ (.D(_00386_),
    .CLK(clknet_leaf_23_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[26][17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11321_ (.D(_00387_),
    .CLK(clknet_leaf_23_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[26][18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11322_ (.D(_00388_),
    .CLK(clknet_leaf_35_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[26][19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11323_ (.D(_00389_),
    .CLK(clknet_leaf_52_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[26][20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11324_ (.D(_00390_),
    .CLK(clknet_leaf_231_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[26][21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11325_ (.D(_00391_),
    .CLK(clknet_leaf_251_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[26][22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11326_ (.D(_00392_),
    .CLK(clknet_leaf_233_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[26][23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11327_ (.D(_00393_),
    .CLK(clknet_leaf_298_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[26][24] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11328_ (.D(_00394_),
    .CLK(clknet_leaf_231_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[26][25] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11329_ (.D(_00395_),
    .CLK(clknet_leaf_292_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[26][26] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11330_ (.D(_00396_),
    .CLK(clknet_leaf_297_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[26][27] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11331_ (.D(_00397_),
    .CLK(clknet_leaf_298_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[26][28] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11332_ (.D(_00398_),
    .CLK(clknet_leaf_186_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[27][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11333_ (.D(_00399_),
    .CLK(clknet_leaf_188_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[27][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11334_ (.D(_00400_),
    .CLK(clknet_leaf_195_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[27][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11335_ (.D(_00401_),
    .CLK(clknet_leaf_140_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[27][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11336_ (.D(_00402_),
    .CLK(clknet_leaf_141_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[27][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11337_ (.D(_00403_),
    .CLK(clknet_leaf_189_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[27][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11338_ (.D(_00404_),
    .CLK(clknet_leaf_201_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[27][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11339_ (.D(_00405_),
    .CLK(clknet_leaf_186_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[27][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11340_ (.D(_00406_),
    .CLK(clknet_leaf_184_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[27][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11341_ (.D(_00407_),
    .CLK(clknet_leaf_199_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[27][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11342_ (.D(_00408_),
    .CLK(clknet_leaf_17_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[27][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11343_ (.D(_00409_),
    .CLK(clknet_leaf_34_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[27][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11344_ (.D(_00410_),
    .CLK(clknet_leaf_0_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[27][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11345_ (.D(_00411_),
    .CLK(clknet_leaf_315_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[27][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11346_ (.D(_00412_),
    .CLK(clknet_leaf_318_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[27][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11347_ (.D(_00413_),
    .CLK(clknet_leaf_313_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[27][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11348_ (.D(_00414_),
    .CLK(clknet_leaf_19_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[27][16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11349_ (.D(_00415_),
    .CLK(clknet_leaf_23_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[27][17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11350_ (.D(_00416_),
    .CLK(clknet_leaf_23_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[27][18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11351_ (.D(_00417_),
    .CLK(clknet_leaf_35_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[27][19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11352_ (.D(_00418_),
    .CLK(clknet_leaf_52_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[27][20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11353_ (.D(_00419_),
    .CLK(clknet_leaf_233_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[27][21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11354_ (.D(_00420_),
    .CLK(clknet_leaf_251_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[27][22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11355_ (.D(_00421_),
    .CLK(clknet_leaf_233_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[27][23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11356_ (.D(_00422_),
    .CLK(clknet_leaf_298_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[27][24] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11357_ (.D(_00423_),
    .CLK(clknet_leaf_231_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[27][25] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11358_ (.D(_00424_),
    .CLK(clknet_leaf_293_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[27][26] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11359_ (.D(_00425_),
    .CLK(clknet_leaf_297_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[27][27] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11360_ (.D(_00426_),
    .CLK(clknet_leaf_298_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[27][28] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11361_ (.D(_00427_),
    .CLK(clknet_leaf_188_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[28][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11362_ (.D(_00428_),
    .CLK(clknet_leaf_224_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[28][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11363_ (.D(_00429_),
    .CLK(clknet_leaf_258_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[28][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11364_ (.D(_00430_),
    .CLK(clknet_leaf_138_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[28][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11365_ (.D(_00431_),
    .CLK(clknet_leaf_195_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[28][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11366_ (.D(_00432_),
    .CLK(clknet_leaf_175_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[28][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11367_ (.D(_00433_),
    .CLK(clknet_leaf_208_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[28][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11368_ (.D(_00434_),
    .CLK(clknet_leaf_186_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[28][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11369_ (.D(_00435_),
    .CLK(clknet_leaf_175_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[28][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11370_ (.D(_00436_),
    .CLK(clknet_leaf_256_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[28][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11371_ (.D(_00437_),
    .CLK(clknet_leaf_12_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[28][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11372_ (.D(_00438_),
    .CLK(clknet_leaf_36_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[28][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11373_ (.D(_00439_),
    .CLK(clknet_leaf_6_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[28][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11374_ (.D(_00440_),
    .CLK(clknet_leaf_311_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[28][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11375_ (.D(_00441_),
    .CLK(clknet_leaf_317_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[28][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11376_ (.D(_00442_),
    .CLK(clknet_leaf_311_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[28][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11377_ (.D(_00443_),
    .CLK(clknet_leaf_30_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[28][16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11378_ (.D(_00444_),
    .CLK(clknet_leaf_73_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[28][17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11379_ (.D(_00445_),
    .CLK(clknet_leaf_30_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[28][18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11380_ (.D(_00446_),
    .CLK(clknet_leaf_71_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[28][19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11381_ (.D(_00447_),
    .CLK(clknet_leaf_52_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[28][20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11382_ (.D(_00448_),
    .CLK(clknet_leaf_291_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[28][21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11383_ (.D(_00449_),
    .CLK(clknet_leaf_270_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[28][22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11384_ (.D(_00450_),
    .CLK(clknet_leaf_290_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[28][23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11385_ (.D(_00451_),
    .CLK(clknet_leaf_300_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[28][24] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11386_ (.D(_00452_),
    .CLK(clknet_leaf_232_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[28][25] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11387_ (.D(_00453_),
    .CLK(clknet_leaf_294_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[28][26] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11388_ (.D(_00454_),
    .CLK(clknet_leaf_272_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[28][27] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11389_ (.D(_00455_),
    .CLK(clknet_leaf_303_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[28][28] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11390_ (.D(_00456_),
    .CLK(clknet_leaf_207_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[2][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11391_ (.D(_00457_),
    .CLK(clknet_leaf_212_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[2][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11392_ (.D(_00458_),
    .CLK(clknet_leaf_258_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[2][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11393_ (.D(_00459_),
    .CLK(clknet_leaf_259_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[2][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11394_ (.D(_00460_),
    .CLK(clknet_leaf_198_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[2][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11395_ (.D(_00461_),
    .CLK(clknet_leaf_212_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[2][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11396_ (.D(_00462_),
    .CLK(clknet_leaf_247_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[2][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11397_ (.D(_00463_),
    .CLK(clknet_leaf_200_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[2][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11398_ (.D(_00464_),
    .CLK(clknet_leaf_220_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[2][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11399_ (.D(_00465_),
    .CLK(clknet_leaf_249_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[2][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11400_ (.D(_00466_),
    .CLK(clknet_leaf_18_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[2][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11401_ (.D(_00467_),
    .CLK(clknet_leaf_14_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[2][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11402_ (.D(_00468_),
    .CLK(clknet_leaf_1_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[2][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11403_ (.D(_00469_),
    .CLK(clknet_leaf_319_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[2][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11404_ (.D(_00470_),
    .CLK(clknet_leaf_320_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[2][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11405_ (.D(_00471_),
    .CLK(clknet_leaf_0_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[2][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11406_ (.D(_00472_),
    .CLK(clknet_leaf_77_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[2][16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11407_ (.D(_00473_),
    .CLK(clknet_leaf_78_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[2][17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11408_ (.D(_00474_),
    .CLK(clknet_leaf_77_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[2][18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11409_ (.D(_00475_),
    .CLK(clknet_leaf_74_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[2][19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11410_ (.D(_00476_),
    .CLK(clknet_leaf_44_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[2][20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11411_ (.D(_00477_),
    .CLK(clknet_leaf_230_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[2][21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11412_ (.D(_00478_),
    .CLK(clknet_leaf_253_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[2][22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11413_ (.D(_00479_),
    .CLK(clknet_leaf_242_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[2][23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11414_ (.D(_00480_),
    .CLK(clknet_leaf_299_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[2][24] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11415_ (.D(_00481_),
    .CLK(clknet_leaf_229_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[2][25] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11416_ (.D(_00482_),
    .CLK(clknet_leaf_295_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[2][26] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11417_ (.D(_00483_),
    .CLK(clknet_leaf_42_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[2][27] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11418_ (.D(_00484_),
    .CLK(clknet_leaf_296_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[2][28] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11419_ (.D(_00485_),
    .CLK(clknet_leaf_187_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[30][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11420_ (.D(_00486_),
    .CLK(clknet_leaf_222_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[30][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11421_ (.D(_00487_),
    .CLK(clknet_leaf_261_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[30][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11422_ (.D(_00488_),
    .CLK(clknet_leaf_135_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[30][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11423_ (.D(_00489_),
    .CLK(clknet_leaf_197_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[30][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11424_ (.D(_00490_),
    .CLK(clknet_leaf_179_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[30][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11425_ (.D(_00491_),
    .CLK(clknet_leaf_210_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[30][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11426_ (.D(_00492_),
    .CLK(clknet_leaf_193_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[30][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11427_ (.D(_00493_),
    .CLK(clknet_leaf_179_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[30][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11428_ (.D(_00494_),
    .CLK(clknet_leaf_255_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[30][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11429_ (.D(_00495_),
    .CLK(clknet_leaf_11_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[30][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11430_ (.D(_00496_),
    .CLK(clknet_leaf_37_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[30][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11431_ (.D(_00497_),
    .CLK(clknet_leaf_6_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[30][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11432_ (.D(_00498_),
    .CLK(clknet_leaf_311_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[30][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11433_ (.D(_00499_),
    .CLK(clknet_leaf_317_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[30][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11434_ (.D(_00500_),
    .CLK(clknet_leaf_309_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[30][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11435_ (.D(_00501_),
    .CLK(clknet_leaf_26_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[30][16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11436_ (.D(_00502_),
    .CLK(clknet_leaf_76_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[30][17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11437_ (.D(_00503_),
    .CLK(clknet_leaf_73_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[30][18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11438_ (.D(_00504_),
    .CLK(clknet_leaf_72_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[30][19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11439_ (.D(_00505_),
    .CLK(clknet_leaf_49_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[30][20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11440_ (.D(_00506_),
    .CLK(clknet_leaf_231_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[30][21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11441_ (.D(_00507_),
    .CLK(clknet_leaf_269_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[30][22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11442_ (.D(_00508_),
    .CLK(clknet_leaf_232_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[30][23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11443_ (.D(_00509_),
    .CLK(clknet_leaf_300_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[30][24] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11444_ (.D(_00510_),
    .CLK(clknet_leaf_231_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[30][25] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11445_ (.D(_00511_),
    .CLK(clknet_leaf_294_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[30][26] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11446_ (.D(_00512_),
    .CLK(clknet_leaf_41_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[30][27] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11447_ (.D(_00513_),
    .CLK(clknet_leaf_302_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[30][28] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11448_ (.D(_00514_),
    .CLK(clknet_leaf_178_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[15][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11449_ (.D(_00515_),
    .CLK(clknet_leaf_222_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[15][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11450_ (.D(_00516_),
    .CLK(clknet_leaf_55_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[15][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11451_ (.D(_00517_),
    .CLK(clknet_leaf_53_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[15][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11452_ (.D(_00518_),
    .CLK(clknet_leaf_53_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[15][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11453_ (.D(_00519_),
    .CLK(clknet_leaf_222_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[15][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11454_ (.D(_00520_),
    .CLK(clknet_leaf_202_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[15][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11455_ (.D(_00521_),
    .CLK(clknet_leaf_192_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[15][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11456_ (.D(_00522_),
    .CLK(clknet_leaf_177_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[15][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11457_ (.D(_00523_),
    .CLK(clknet_leaf_257_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[15][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11458_ (.D(_00524_),
    .CLK(clknet_leaf_15_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[15][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11459_ (.D(_00525_),
    .CLK(clknet_leaf_33_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[15][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11460_ (.D(_00526_),
    .CLK(clknet_leaf_308_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[15][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11461_ (.D(_00527_),
    .CLK(clknet_leaf_10_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[15][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11462_ (.D(_00528_),
    .CLK(clknet_leaf_309_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[15][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11463_ (.D(_00529_),
    .CLK(clknet_leaf_9_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[15][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11464_ (.D(_00530_),
    .CLK(clknet_leaf_20_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[15][16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11465_ (.D(_00531_),
    .CLK(clknet_leaf_20_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[15][17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11466_ (.D(_00532_),
    .CLK(clknet_leaf_22_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[15][18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11467_ (.D(_00533_),
    .CLK(clknet_leaf_29_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[15][19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11468_ (.D(_00534_),
    .CLK(clknet_leaf_50_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[15][20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11469_ (.D(_00535_),
    .CLK(clknet_leaf_283_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[15][21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11470_ (.D(_00536_),
    .CLK(clknet_leaf_268_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[15][22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11471_ (.D(_00537_),
    .CLK(clknet_leaf_284_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[15][23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11472_ (.D(_00538_),
    .CLK(clknet_leaf_305_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[15][24] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11473_ (.D(_00539_),
    .CLK(clknet_leaf_285_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[15][25] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11474_ (.D(_00540_),
    .CLK(clknet_leaf_281_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[15][26] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11475_ (.D(_00541_),
    .CLK(clknet_leaf_42_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[15][27] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11476_ (.D(_00542_),
    .CLK(clknet_leaf_270_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[15][28] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11477_ (.D(_00543_),
    .CLK(clknet_leaf_187_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[24][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11478_ (.D(_00544_),
    .CLK(clknet_leaf_180_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[24][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11479_ (.D(_00545_),
    .CLK(clknet_leaf_196_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[24][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11480_ (.D(_00546_),
    .CLK(clknet_leaf_141_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[24][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11481_ (.D(_00547_),
    .CLK(clknet_leaf_141_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[24][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11482_ (.D(_00548_),
    .CLK(clknet_leaf_179_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[24][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11483_ (.D(_00549_),
    .CLK(clknet_leaf_201_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[24][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11484_ (.D(_00550_),
    .CLK(clknet_leaf_185_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[24][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11485_ (.D(_00551_),
    .CLK(clknet_leaf_180_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[24][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11486_ (.D(_00552_),
    .CLK(clknet_leaf_201_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[24][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11487_ (.D(_00553_),
    .CLK(clknet_leaf_17_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[24][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11488_ (.D(_00554_),
    .CLK(clknet_leaf_33_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[24][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11489_ (.D(_00555_),
    .CLK(clknet_leaf_319_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[24][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11490_ (.D(_00556_),
    .CLK(clknet_leaf_314_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[24][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11491_ (.D(_00557_),
    .CLK(clknet_leaf_318_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[24][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11492_ (.D(_00558_),
    .CLK(clknet_leaf_313_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[24][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11493_ (.D(_00559_),
    .CLK(clknet_leaf_20_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[24][16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11494_ (.D(_00560_),
    .CLK(clknet_leaf_19_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[24][17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11495_ (.D(_00561_),
    .CLK(clknet_leaf_23_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[24][18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11496_ (.D(_00562_),
    .CLK(clknet_leaf_34_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[24][19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11497_ (.D(_00563_),
    .CLK(clknet_leaf_261_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[24][20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11498_ (.D(_00564_),
    .CLK(clknet_leaf_230_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[24][21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11499_ (.D(_00565_),
    .CLK(clknet_leaf_251_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[24][22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11500_ (.D(_00566_),
    .CLK(clknet_leaf_234_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[24][23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11501_ (.D(_00567_),
    .CLK(clknet_leaf_298_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[24][24] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11502_ (.D(_00568_),
    .CLK(clknet_leaf_230_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[24][25] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11503_ (.D(_00569_),
    .CLK(clknet_leaf_292_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[24][26] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11504_ (.D(_00570_),
    .CLK(clknet_leaf_293_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[24][27] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11505_ (.D(_00571_),
    .CLK(clknet_leaf_297_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[24][28] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11506_ (.D(_00572_),
    .CLK(clknet_5_22_0_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[23][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11507_ (.D(_00573_),
    .CLK(clknet_leaf_211_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[23][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11508_ (.D(_00574_),
    .CLK(clknet_leaf_55_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[23][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11509_ (.D(_00575_),
    .CLK(clknet_leaf_134_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[23][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11510_ (.D(_00576_),
    .CLK(clknet_leaf_134_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[23][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11511_ (.D(_00577_),
    .CLK(clknet_leaf_213_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[23][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11512_ (.D(_00578_),
    .CLK(clknet_leaf_247_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[23][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11513_ (.D(_00579_),
    .CLK(clknet_leaf_195_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[23][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11514_ (.D(_00580_),
    .CLK(clknet_leaf_208_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[23][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11515_ (.D(_00581_),
    .CLK(clknet_leaf_253_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[23][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11516_ (.D(_00582_),
    .CLK(clknet_leaf_14_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[23][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11517_ (.D(_00583_),
    .CLK(clknet_leaf_37_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[23][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11518_ (.D(_00584_),
    .CLK(clknet_leaf_306_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[23][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11519_ (.D(_00585_),
    .CLK(clknet_leaf_39_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[23][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11520_ (.D(_00586_),
    .CLK(clknet_leaf_3_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[23][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11521_ (.D(_00587_),
    .CLK(clknet_leaf_307_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[23][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11522_ (.D(_00588_),
    .CLK(clknet_leaf_29_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[23][16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11523_ (.D(_00589_),
    .CLK(clknet_leaf_29_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[23][17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11524_ (.D(_00590_),
    .CLK(clknet_leaf_27_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[23][18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11525_ (.D(_00591_),
    .CLK(clknet_leaf_32_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[23][19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11526_ (.D(_00592_),
    .CLK(clknet_leaf_50_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[23][20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11527_ (.D(_00593_),
    .CLK(clknet_leaf_240_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[23][21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11528_ (.D(_00594_),
    .CLK(clknet_leaf_240_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[23][22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11529_ (.D(_00595_),
    .CLK(clknet_leaf_243_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[23][23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11530_ (.D(_00596_),
    .CLK(clknet_leaf_278_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[23][24] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11531_ (.D(_00597_),
    .CLK(clknet_leaf_242_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[23][25] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11532_ (.D(_00598_),
    .CLK(clknet_leaf_281_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[23][26] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11533_ (.D(_00599_),
    .CLK(clknet_leaf_272_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[23][27] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11534_ (.D(_00600_),
    .CLK(clknet_leaf_277_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[23][28] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11535_ (.D(_00601_),
    .CLK(clknet_leaf_184_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[25][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11536_ (.D(_00602_),
    .CLK(clknet_leaf_180_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[25][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11537_ (.D(_00603_),
    .CLK(clknet_leaf_196_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[25][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11538_ (.D(_00604_),
    .CLK(clknet_leaf_142_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[25][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11539_ (.D(_00605_),
    .CLK(clknet_leaf_141_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[25][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11540_ (.D(_00606_),
    .CLK(clknet_leaf_179_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[25][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11541_ (.D(_00607_),
    .CLK(clknet_leaf_201_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[25][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11542_ (.D(_00608_),
    .CLK(clknet_leaf_146_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[25][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11543_ (.D(_00609_),
    .CLK(clknet_5_29_0_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[25][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11544_ (.D(_00610_),
    .CLK(clknet_leaf_257_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[25][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11545_ (.D(_00611_),
    .CLK(clknet_leaf_17_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[25][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11546_ (.D(_00612_),
    .CLK(clknet_leaf_33_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[25][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11547_ (.D(_00613_),
    .CLK(clknet_leaf_319_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[25][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11548_ (.D(_00614_),
    .CLK(clknet_leaf_315_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[25][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11549_ (.D(_00615_),
    .CLK(clknet_leaf_318_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[25][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11550_ (.D(_00616_),
    .CLK(clknet_leaf_313_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[25][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11551_ (.D(_00617_),
    .CLK(clknet_leaf_18_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[25][16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11552_ (.D(_00618_),
    .CLK(clknet_leaf_22_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[25][17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11553_ (.D(_00619_),
    .CLK(clknet_leaf_23_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[25][18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11554_ (.D(_00620_),
    .CLK(clknet_leaf_35_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[25][19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11555_ (.D(_00621_),
    .CLK(clknet_leaf_263_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[25][20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11556_ (.D(_00622_),
    .CLK(clknet_leaf_230_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[25][21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11557_ (.D(_00623_),
    .CLK(clknet_leaf_251_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[25][22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11558_ (.D(_00624_),
    .CLK(clknet_leaf_233_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[25][23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11559_ (.D(_00625_),
    .CLK(clknet_leaf_298_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[25][24] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11560_ (.D(_00626_),
    .CLK(clknet_leaf_231_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[25][25] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11561_ (.D(_00627_),
    .CLK(clknet_leaf_292_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[25][26] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11562_ (.D(_00628_),
    .CLK(clknet_leaf_293_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[25][27] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11563_ (.D(_00629_),
    .CLK(clknet_leaf_297_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[25][28] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11564_ (.D(_00630_),
    .CLK(clknet_leaf_205_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[22][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11565_ (.D(_00631_),
    .CLK(clknet_leaf_208_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[22][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11566_ (.D(_00632_),
    .CLK(clknet_leaf_55_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[22][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11567_ (.D(_00633_),
    .CLK(clknet_leaf_134_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[22][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11568_ (.D(_00634_),
    .CLK(clknet_leaf_134_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[22][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11569_ (.D(_00635_),
    .CLK(clknet_leaf_211_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[22][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11570_ (.D(_00636_),
    .CLK(clknet_leaf_248_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[22][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11571_ (.D(_00637_),
    .CLK(clknet_leaf_194_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[22][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11572_ (.D(_00638_),
    .CLK(clknet_leaf_208_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[22][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11573_ (.D(_00639_),
    .CLK(clknet_leaf_254_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[22][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11574_ (.D(_00640_),
    .CLK(clknet_leaf_20_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[22][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11575_ (.D(_00641_),
    .CLK(clknet_leaf_34_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[22][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11576_ (.D(_00642_),
    .CLK(clknet_leaf_307_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[22][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11577_ (.D(_00643_),
    .CLK(clknet_leaf_40_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[22][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11578_ (.D(_00644_),
    .CLK(clknet_leaf_8_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[22][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11579_ (.D(_00645_),
    .CLK(clknet_leaf_276_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[22][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11580_ (.D(_00646_),
    .CLK(clknet_leaf_26_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[22][16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11581_ (.D(_00647_),
    .CLK(clknet_leaf_26_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[22][17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11582_ (.D(_00648_),
    .CLK(clknet_leaf_27_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[22][18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11583_ (.D(_00649_),
    .CLK(clknet_leaf_29_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[22][19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11584_ (.D(_00650_),
    .CLK(clknet_leaf_50_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[22][20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11585_ (.D(_00651_),
    .CLK(clknet_leaf_240_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[22][21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11586_ (.D(_00652_),
    .CLK(clknet_leaf_240_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[22][22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11587_ (.D(_00653_),
    .CLK(clknet_leaf_241_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[22][23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11588_ (.D(_00654_),
    .CLK(clknet_leaf_277_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[22][24] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11589_ (.D(_00655_),
    .CLK(clknet_leaf_242_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[22][25] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11590_ (.D(_00656_),
    .CLK(clknet_leaf_281_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[22][26] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11591_ (.D(_00657_),
    .CLK(clknet_leaf_44_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[22][27] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11592_ (.D(_00658_),
    .CLK(clknet_leaf_276_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[22][28] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11593_ (.D(_00659_),
    .CLK(clknet_leaf_205_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[21][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11594_ (.D(_00660_),
    .CLK(clknet_leaf_208_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[21][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11595_ (.D(_00661_),
    .CLK(clknet_leaf_136_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[21][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11596_ (.D(_00662_),
    .CLK(clknet_leaf_132_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[21][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11597_ (.D(_00663_),
    .CLK(clknet_leaf_132_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[21][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11598_ (.D(_00664_),
    .CLK(clknet_leaf_212_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[21][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11599_ (.D(_00665_),
    .CLK(clknet_leaf_248_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[21][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11600_ (.D(_00666_),
    .CLK(clknet_leaf_194_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[21][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11601_ (.D(_00667_),
    .CLK(clknet_leaf_207_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[21][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11602_ (.D(_00668_),
    .CLK(clknet_leaf_254_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[21][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11603_ (.D(_00669_),
    .CLK(clknet_leaf_20_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[21][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11604_ (.D(_00670_),
    .CLK(clknet_leaf_34_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[21][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11605_ (.D(_00671_),
    .CLK(clknet_leaf_306_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[21][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11606_ (.D(_00672_),
    .CLK(clknet_leaf_41_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[21][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11607_ (.D(_00673_),
    .CLK(clknet_leaf_308_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[21][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11608_ (.D(_00674_),
    .CLK(clknet_leaf_307_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[21][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11609_ (.D(_00675_),
    .CLK(clknet_leaf_26_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[21][16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11610_ (.D(_00676_),
    .CLK(clknet_leaf_27_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[21][17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11611_ (.D(_00677_),
    .CLK(clknet_leaf_28_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[21][18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11612_ (.D(_00678_),
    .CLK(clknet_leaf_31_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[21][19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11613_ (.D(_00679_),
    .CLK(clknet_leaf_50_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[21][20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11614_ (.D(_00680_),
    .CLK(clknet_leaf_239_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[21][21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11615_ (.D(_00681_),
    .CLK(clknet_leaf_250_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[21][22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11616_ (.D(_00682_),
    .CLK(clknet_leaf_241_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[21][23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11617_ (.D(_00683_),
    .CLK(clknet_leaf_303_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[21][24] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11618_ (.D(_00684_),
    .CLK(clknet_leaf_241_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[21][25] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11619_ (.D(_00685_),
    .CLK(clknet_leaf_287_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[21][26] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11620_ (.D(_00686_),
    .CLK(clknet_leaf_44_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[21][27] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11621_ (.D(_00687_),
    .CLK(clknet_leaf_274_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[21][28] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11622_ (.D(_00688_),
    .CLK(clknet_leaf_47_wb_clk_i),
    .Q(_00000_));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11623_ (.D(_00689_),
    .CLK(clknet_leaf_47_wb_clk_i),
    .Q(_00001_));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11624_ (.D(_00690_),
    .CLK(clknet_leaf_32_wb_clk_i),
    .Q(_00002_));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11625_ (.D(_00691_),
    .CLK(clknet_leaf_32_wb_clk_i),
    .Q(_00003_));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11626_ (.D(_00692_),
    .CLK(clknet_leaf_32_wb_clk_i),
    .Q(_00004_));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11627_ (.D(_00005_),
    .CLK(clknet_leaf_62_wb_clk_i),
    .Q(\soc.spi_video_ram_1.current_state[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11628_ (.D(_00006_),
    .CLK(clknet_leaf_62_wb_clk_i),
    .Q(\soc.spi_video_ram_1.current_state[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11629_ (.D(_00007_),
    .CLK(clknet_leaf_69_wb_clk_i),
    .Q(\soc.spi_video_ram_1.current_state[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11630_ (.D(_00008_),
    .CLK(clknet_leaf_64_wb_clk_i),
    .Q(\soc.spi_video_ram_1.current_state[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11631_ (.D(_00009_),
    .CLK(clknet_leaf_62_wb_clk_i),
    .Q(\soc.spi_video_ram_1.current_state[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11632_ (.D(_00693_),
    .CLK(clknet_leaf_207_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[20][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11633_ (.D(_00694_),
    .CLK(clknet_leaf_216_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[20][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11634_ (.D(_00695_),
    .CLK(clknet_leaf_137_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[20][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11635_ (.D(_00696_),
    .CLK(clknet_leaf_139_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[20][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11636_ (.D(_00697_),
    .CLK(clknet_leaf_139_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[20][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11637_ (.D(_00698_),
    .CLK(clknet_leaf_215_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[20][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11638_ (.D(_00699_),
    .CLK(clknet_leaf_210_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[20][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11639_ (.D(_00700_),
    .CLK(clknet_leaf_195_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[20][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11640_ (.D(_00701_),
    .CLK(clknet_leaf_208_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[20][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11641_ (.D(_00702_),
    .CLK(clknet_leaf_256_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[20][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11642_ (.D(_00703_),
    .CLK(clknet_leaf_14_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[20][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11643_ (.D(_00704_),
    .CLK(clknet_leaf_36_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[20][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11644_ (.D(_00705_),
    .CLK(clknet_leaf_308_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[20][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11645_ (.D(_00706_),
    .CLK(clknet_leaf_39_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[20][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11646_ (.D(_00707_),
    .CLK(clknet_leaf_6_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[20][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11647_ (.D(_00708_),
    .CLK(clknet_leaf_308_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[20][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11648_ (.D(_00709_),
    .CLK(clknet_leaf_29_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[20][16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11649_ (.D(_00710_),
    .CLK(clknet_leaf_27_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[20][17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11650_ (.D(_00711_),
    .CLK(clknet_leaf_28_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[20][18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11651_ (.D(_00712_),
    .CLK(clknet_leaf_32_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[20][19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11652_ (.D(_00713_),
    .CLK(clknet_leaf_51_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[20][20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11653_ (.D(_00714_),
    .CLK(clknet_leaf_239_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[20][21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11654_ (.D(_00715_),
    .CLK(clknet_leaf_249_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[20][22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11655_ (.D(_00716_),
    .CLK(clknet_leaf_239_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[20][23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11656_ (.D(_00717_),
    .CLK(clknet_leaf_304_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[20][24] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11657_ (.D(_00718_),
    .CLK(clknet_leaf_235_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[20][25] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11658_ (.D(_00719_),
    .CLK(clknet_leaf_287_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[20][26] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11659_ (.D(_00720_),
    .CLK(clknet_leaf_272_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[20][27] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11660_ (.D(_00721_),
    .CLK(clknet_leaf_276_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[20][28] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11661_ (.D(_00722_),
    .CLK(clknet_leaf_65_wb_clk_i),
    .Q(\soc.spi_video_ram_1.state_counter[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11662_ (.D(_00723_),
    .CLK(clknet_leaf_64_wb_clk_i),
    .Q(\soc.spi_video_ram_1.state_counter[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11663_ (.D(_00724_),
    .CLK(clknet_leaf_65_wb_clk_i),
    .Q(\soc.spi_video_ram_1.state_counter[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11664_ (.D(_00725_),
    .CLK(clknet_leaf_66_wb_clk_i),
    .Q(\soc.spi_video_ram_1.state_counter[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11665_ (.D(_00726_),
    .CLK(clknet_leaf_67_wb_clk_i),
    .Q(\soc.spi_video_ram_1.state_counter[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11666_ (.D(_00727_),
    .CLK(clknet_leaf_83_wb_clk_i),
    .Q(\soc.spi_video_ram_1.state_counter[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11667_ (.D(_00728_),
    .CLK(clknet_leaf_66_wb_clk_i),
    .Q(\soc.spi_video_ram_1.state_counter[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11668_ (.D(_00729_),
    .CLK(clknet_leaf_66_wb_clk_i),
    .Q(\soc.spi_video_ram_1.state_counter[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11669_ (.D(_00730_),
    .CLK(clknet_leaf_64_wb_clk_i),
    .Q(\soc.spi_video_ram_1.state_counter[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11670_ (.D(_00731_),
    .CLK(clknet_leaf_65_wb_clk_i),
    .Q(\soc.spi_video_ram_1.state_counter[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11671_ (.D(_00732_),
    .CLK(clknet_leaf_66_wb_clk_i),
    .Q(\soc.spi_video_ram_1.state_counter[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11672_ (.D(_00733_),
    .CLK(clknet_leaf_127_wb_clk_i),
    .Q(\soc.video_generator_1.v_count[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11673_ (.D(_00734_),
    .CLK(clknet_leaf_128_wb_clk_i),
    .Q(\soc.video_generator_1.v_count[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11674_ (.D(_00735_),
    .CLK(clknet_leaf_128_wb_clk_i),
    .Q(\soc.video_generator_1.v_count[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11675_ (.D(_00736_),
    .CLK(clknet_leaf_129_wb_clk_i),
    .Q(\soc.video_generator_1.v_count[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11676_ (.D(_00737_),
    .CLK(clknet_leaf_64_wb_clk_i),
    .Q(\soc.video_generator_1.v_count[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11677_ (.D(_00738_),
    .CLK(clknet_leaf_64_wb_clk_i),
    .Q(\soc.video_generator_1.v_count[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11678_ (.D(_00739_),
    .CLK(clknet_leaf_64_wb_clk_i),
    .Q(\soc.video_generator_1.v_count[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11679_ (.D(_00740_),
    .CLK(clknet_leaf_63_wb_clk_i),
    .Q(\soc.video_generator_1.v_count[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11680_ (.D(_00741_),
    .CLK(clknet_leaf_63_wb_clk_i),
    .Q(\soc.video_generator_1.v_count[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11681_ (.D(_00742_),
    .CLK(clknet_leaf_129_wb_clk_i),
    .Q(\soc.video_generator_1.v_count[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11682_ (.D(_00743_),
    .CLK(clknet_leaf_186_wb_clk_i),
    .Q(\soc.spi_video_ram_1.fifo_in_data[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11683_ (.D(_00744_),
    .CLK(clknet_leaf_145_wb_clk_i),
    .Q(\soc.spi_video_ram_1.fifo_in_data[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11684_ (.D(_00745_),
    .CLK(clknet_leaf_143_wb_clk_i),
    .Q(\soc.spi_video_ram_1.fifo_in_data[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11685_ (.D(_00746_),
    .CLK(clknet_leaf_132_wb_clk_i),
    .Q(\soc.spi_video_ram_1.fifo_in_data[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11686_ (.D(_00747_),
    .CLK(clknet_leaf_142_wb_clk_i),
    .Q(\soc.spi_video_ram_1.fifo_in_data[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11687_ (.D(_00748_),
    .CLK(clknet_leaf_146_wb_clk_i),
    .Q(\soc.spi_video_ram_1.fifo_in_data[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11688_ (.D(_00749_),
    .CLK(clknet_leaf_145_wb_clk_i),
    .Q(\soc.spi_video_ram_1.fifo_in_data[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11689_ (.D(_00750_),
    .CLK(clknet_leaf_145_wb_clk_i),
    .Q(\soc.spi_video_ram_1.fifo_in_data[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11690_ (.D(_00751_),
    .CLK(clknet_leaf_145_wb_clk_i),
    .Q(\soc.spi_video_ram_1.fifo_in_data[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11691_ (.D(_00752_),
    .CLK(clknet_leaf_141_wb_clk_i),
    .Q(\soc.spi_video_ram_1.fifo_in_data[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11692_ (.D(_00753_),
    .CLK(clknet_leaf_132_wb_clk_i),
    .Q(\soc.spi_video_ram_1.fifo_in_data[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11693_ (.D(_00754_),
    .CLK(clknet_leaf_130_wb_clk_i),
    .Q(\soc.spi_video_ram_1.fifo_in_data[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11694_ (.D(_00755_),
    .CLK(clknet_leaf_304_wb_clk_i),
    .Q(\soc.spi_video_ram_1.fifo_in_data[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11695_ (.D(_00756_),
    .CLK(clknet_leaf_301_wb_clk_i),
    .Q(\soc.spi_video_ram_1.fifo_in_data[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11696_ (.D(_00757_),
    .CLK(clknet_leaf_300_wb_clk_i),
    .Q(\soc.spi_video_ram_1.fifo_in_data[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11697_ (.D(_00758_),
    .CLK(clknet_leaf_300_wb_clk_i),
    .Q(\soc.spi_video_ram_1.fifo_in_data[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11698_ (.D(_00759_),
    .CLK(clknet_leaf_191_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[9][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11699_ (.D(_00760_),
    .CLK(clknet_5_22_0_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[9][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11700_ (.D(_00761_),
    .CLK(clknet_leaf_198_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[9][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11701_ (.D(_00762_),
    .CLK(clknet_leaf_198_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[9][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11702_ (.D(_00763_),
    .CLK(clknet_leaf_200_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[9][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11703_ (.D(_00764_),
    .CLK(clknet_leaf_222_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[9][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11704_ (.D(_00765_),
    .CLK(clknet_leaf_205_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[9][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11705_ (.D(_00766_),
    .CLK(clknet_leaf_191_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[9][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11706_ (.D(_00767_),
    .CLK(clknet_leaf_178_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[9][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11707_ (.D(_00768_),
    .CLK(clknet_leaf_256_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[9][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11708_ (.D(_00769_),
    .CLK(clknet_leaf_17_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[9][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11709_ (.D(_00770_),
    .CLK(clknet_leaf_42_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[9][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11710_ (.D(_00771_),
    .CLK(clknet_leaf_2_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[9][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11711_ (.D(_00772_),
    .CLK(clknet_leaf_8_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[9][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11712_ (.D(_00773_),
    .CLK(clknet_leaf_7_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[9][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11713_ (.D(_00774_),
    .CLK(clknet_leaf_9_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[9][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11714_ (.D(_00775_),
    .CLK(clknet_leaf_76_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[9][16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11715_ (.D(_00776_),
    .CLK(clknet_leaf_24_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[9][17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11716_ (.D(_00777_),
    .CLK(clknet_leaf_25_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[9][18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11717_ (.D(_00778_),
    .CLK(clknet_leaf_32_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[9][19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11718_ (.D(_00779_),
    .CLK(clknet_leaf_53_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[9][20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11719_ (.D(_00780_),
    .CLK(clknet_leaf_283_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[9][21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11720_ (.D(_00781_),
    .CLK(clknet_leaf_238_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[9][22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11721_ (.D(_00782_),
    .CLK(clknet_leaf_238_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[9][23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11722_ (.D(_00783_),
    .CLK(clknet_leaf_276_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[9][24] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11723_ (.D(_00784_),
    .CLK(clknet_leaf_239_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[9][25] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11724_ (.D(_00785_),
    .CLK(clknet_leaf_281_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[9][26] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11725_ (.D(_00786_),
    .CLK(clknet_leaf_272_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[9][27] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11726_ (.D(_00787_),
    .CLK(clknet_leaf_274_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[9][28] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11727_ (.D(_00788_),
    .CLK(clknet_leaf_214_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[4][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11728_ (.D(_00789_),
    .CLK(clknet_leaf_227_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[4][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11729_ (.D(_00790_),
    .CLK(clknet_leaf_254_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[4][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11730_ (.D(_00791_),
    .CLK(clknet_leaf_262_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[4][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11731_ (.D(_00792_),
    .CLK(clknet_leaf_262_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[4][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11732_ (.D(_00793_),
    .CLK(clknet_leaf_227_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[4][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11733_ (.D(_00794_),
    .CLK(clknet_leaf_245_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[4][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11734_ (.D(_00795_),
    .CLK(clknet_leaf_244_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[4][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11735_ (.D(_00796_),
    .CLK(clknet_leaf_228_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[4][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11736_ (.D(_00797_),
    .CLK(clknet_leaf_246_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[4][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11737_ (.D(_00798_),
    .CLK(clknet_leaf_15_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[4][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11738_ (.D(_00799_),
    .CLK(clknet_leaf_39_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[4][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11739_ (.D(_00800_),
    .CLK(clknet_leaf_308_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[4][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11740_ (.D(_00801_),
    .CLK(clknet_leaf_314_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[4][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11741_ (.D(_00802_),
    .CLK(clknet_leaf_315_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[4][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11742_ (.D(_00803_),
    .CLK(clknet_leaf_316_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[4][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11743_ (.D(_00804_),
    .CLK(clknet_leaf_74_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[4][16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11744_ (.D(_00805_),
    .CLK(clknet_leaf_67_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[4][17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11745_ (.D(_00806_),
    .CLK(clknet_leaf_75_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[4][18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11746_ (.D(_00807_),
    .CLK(clknet_leaf_70_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[4][19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11747_ (.D(_00808_),
    .CLK(clknet_leaf_59_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[4][20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11748_ (.D(_00809_),
    .CLK(clknet_leaf_289_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[4][21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11749_ (.D(_00810_),
    .CLK(clknet_leaf_267_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[4][22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11750_ (.D(_00811_),
    .CLK(clknet_leaf_287_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[4][23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11751_ (.D(_00812_),
    .CLK(clknet_leaf_302_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[4][24] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11752_ (.D(_00813_),
    .CLK(clknet_leaf_287_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[4][25] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11753_ (.D(_00814_),
    .CLK(clknet_leaf_295_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[4][26] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11754_ (.D(_00815_),
    .CLK(clknet_5_6_0_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[4][27] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11755_ (.D(_00816_),
    .CLK(clknet_leaf_279_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[4][28] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11756_ (.D(_00817_),
    .CLK(clknet_leaf_100_wb_clk_i),
    .Q(\soc.rom_loader.was_loading ));
 gf180mcu_fd_sc_mcu7t5v0__dffnq_2 _11757_ (.D(_00818_),
    .CLKN(clknet_leaf_61_wb_clk_i),
    .Q(\soc.spi_video_ram_1.state_sram_clk_counter[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffnq_2 _11758_ (.D(_00819_),
    .CLKN(clknet_leaf_61_wb_clk_i),
    .Q(\soc.spi_video_ram_1.state_sram_clk_counter[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffnq_1 _11759_ (.D(_00820_),
    .CLKN(clknet_leaf_71_wb_clk_i),
    .Q(\soc.spi_video_ram_1.state_sram_clk_counter[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffnq_2 _11760_ (.D(_00821_),
    .CLKN(clknet_leaf_70_wb_clk_i),
    .Q(\soc.spi_video_ram_1.state_sram_clk_counter[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffnq_1 _11761_ (.D(_00822_),
    .CLKN(clknet_leaf_70_wb_clk_i),
    .Q(\soc.spi_video_ram_1.state_sram_clk_counter[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffnq_1 _11762_ (.D(_00823_),
    .CLKN(clknet_leaf_70_wb_clk_i),
    .Q(\soc.spi_video_ram_1.state_sram_clk_counter[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffnq_1 _11763_ (.D(_00824_),
    .CLKN(clknet_leaf_68_wb_clk_i),
    .Q(\soc.spi_video_ram_1.state_sram_clk_counter[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffnq_2 _11764_ (.D(_00825_),
    .CLKN(clknet_leaf_68_wb_clk_i),
    .Q(\soc.spi_video_ram_1.state_sram_clk_counter[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffnq_1 _11765_ (.D(_00826_),
    .CLKN(clknet_leaf_69_wb_clk_i),
    .Q(\soc.spi_video_ram_1.state_sram_clk_counter[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffnq_1 _11766_ (.D(_00827_),
    .CLKN(clknet_leaf_69_wb_clk_i),
    .Q(net69));
 gf180mcu_fd_sc_mcu7t5v0__dffnq_1 _11767_ (.D(_00828_),
    .CLKN(clknet_leaf_63_wb_clk_i),
    .Q(\soc.spi_video_ram_1.sram_sck_rise_edge ));
 gf180mcu_fd_sc_mcu7t5v0__dffnq_1 _11768_ (.D(_00829_),
    .CLKN(clknet_leaf_69_wb_clk_i),
    .Q(\soc.spi_video_ram_1.sram_sck_fall_edge ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11769_ (.D(_00830_),
    .CLK(clknet_leaf_60_wb_clk_i),
    .Q(net68));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11770_ (.D(_00831_),
    .CLK(clknet_leaf_89_wb_clk_i),
    .Q(\soc.spi_video_ram_1.read_value[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11771_ (.D(_00832_),
    .CLK(clknet_leaf_82_wb_clk_i),
    .Q(\soc.spi_video_ram_1.read_value[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11772_ (.D(_00833_),
    .CLK(clknet_leaf_81_wb_clk_i),
    .Q(\soc.spi_video_ram_1.read_value[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11773_ (.D(_00834_),
    .CLK(clknet_leaf_89_wb_clk_i),
    .Q(\soc.spi_video_ram_1.read_value[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11774_ (.D(_00835_),
    .CLK(clknet_leaf_105_wb_clk_i),
    .Q(\soc.rom_encoder_0.output_buffer[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11775_ (.D(_00836_),
    .CLK(clknet_leaf_107_wb_clk_i),
    .Q(\soc.rom_encoder_0.output_buffer[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11776_ (.D(_00837_),
    .CLK(clknet_leaf_93_wb_clk_i),
    .Q(\soc.rom_encoder_0.output_buffer[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11777_ (.D(_00838_),
    .CLK(clknet_leaf_104_wb_clk_i),
    .Q(\soc.rom_encoder_0.output_buffer[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11778_ (.D(_00839_),
    .CLK(clknet_leaf_93_wb_clk_i),
    .Q(\soc.rom_encoder_0.output_buffer[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11779_ (.D(_00840_),
    .CLK(clknet_leaf_104_wb_clk_i),
    .Q(\soc.rom_encoder_0.output_buffer[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11780_ (.D(_00841_),
    .CLK(clknet_leaf_104_wb_clk_i),
    .Q(\soc.rom_encoder_0.output_buffer[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11781_ (.D(_00842_),
    .CLK(clknet_leaf_104_wb_clk_i),
    .Q(\soc.rom_encoder_0.output_buffer[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11782_ (.D(_00843_),
    .CLK(clknet_5_14_0_wb_clk_i),
    .Q(\soc.rom_encoder_0.output_buffer[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11783_ (.D(_00844_),
    .CLK(clknet_leaf_104_wb_clk_i),
    .Q(\soc.rom_encoder_0.output_buffer[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11784_ (.D(_00845_),
    .CLK(clknet_leaf_102_wb_clk_i),
    .Q(\soc.rom_encoder_0.output_buffer[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11785_ (.D(_00846_),
    .CLK(clknet_leaf_98_wb_clk_i),
    .Q(\soc.rom_encoder_0.output_buffer[16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11786_ (.D(_00847_),
    .CLK(clknet_leaf_104_wb_clk_i),
    .Q(\soc.rom_encoder_0.output_buffer[17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11787_ (.D(_00848_),
    .CLK(clknet_leaf_102_wb_clk_i),
    .Q(\soc.rom_encoder_0.output_buffer[18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11788_ (.D(_00849_),
    .CLK(clknet_leaf_101_wb_clk_i),
    .Q(\soc.rom_encoder_0.output_buffer[19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11789_ (.D(_00850_),
    .CLK(clknet_leaf_63_wb_clk_i),
    .Q(\soc.spi_video_ram_1.buffer_index[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11790_ (.D(_00851_),
    .CLK(clknet_leaf_63_wb_clk_i),
    .Q(\soc.spi_video_ram_1.buffer_index[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11791_ (.D(_00852_),
    .CLK(clknet_leaf_130_wb_clk_i),
    .Q(\soc.spi_video_ram_1.buffer_index[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11792_ (.D(_00853_),
    .CLK(clknet_leaf_130_wb_clk_i),
    .Q(\soc.spi_video_ram_1.buffer_index[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11793_ (.D(_00854_),
    .CLK(clknet_leaf_130_wb_clk_i),
    .Q(\soc.spi_video_ram_1.buffer_index[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11794_ (.D(_00855_),
    .CLK(clknet_5_24_0_wb_clk_i),
    .Q(\soc.spi_video_ram_1.buffer_index[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11795_ (.D(_00011_),
    .CLK(clknet_leaf_132_wb_clk_i),
    .Q(\soc.spi_video_ram_1.fifo_write_request ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11796_ (.D(_00856_),
    .CLK(clknet_leaf_71_wb_clk_i),
    .Q(\soc.spi_video_ram_1.sram_sio_oe ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11797_ (.D(_00857_),
    .CLK(clknet_leaf_82_wb_clk_i),
    .Q(\soc.spi_video_ram_1.fifo_in_address[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11798_ (.D(_00858_),
    .CLK(clknet_leaf_83_wb_clk_i),
    .Q(\soc.spi_video_ram_1.fifo_in_address[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11799_ (.D(_00859_),
    .CLK(clknet_leaf_74_wb_clk_i),
    .Q(\soc.spi_video_ram_1.fifo_in_address[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11800_ (.D(_00860_),
    .CLK(clknet_leaf_67_wb_clk_i),
    .Q(\soc.spi_video_ram_1.fifo_in_address[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11801_ (.D(_00861_),
    .CLK(clknet_leaf_55_wb_clk_i),
    .Q(\soc.spi_video_ram_1.fifo_in_address[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11802_ (.D(_00862_),
    .CLK(clknet_leaf_291_wb_clk_i),
    .Q(\soc.spi_video_ram_1.fifo_in_address[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11803_ (.D(_00863_),
    .CLK(clknet_leaf_265_wb_clk_i),
    .Q(\soc.spi_video_ram_1.fifo_in_address[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11804_ (.D(_00864_),
    .CLK(clknet_leaf_286_wb_clk_i),
    .Q(\soc.spi_video_ram_1.fifo_in_address[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11805_ (.D(_00865_),
    .CLK(clknet_leaf_295_wb_clk_i),
    .Q(\soc.spi_video_ram_1.fifo_in_address[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11806_ (.D(_00866_),
    .CLK(clknet_leaf_288_wb_clk_i),
    .Q(\soc.spi_video_ram_1.fifo_in_address[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11807_ (.D(_00867_),
    .CLK(clknet_leaf_288_wb_clk_i),
    .Q(\soc.spi_video_ram_1.fifo_in_address[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11808_ (.D(_00868_),
    .CLK(clknet_leaf_263_wb_clk_i),
    .Q(\soc.spi_video_ram_1.fifo_in_address[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11809_ (.D(_00869_),
    .CLK(clknet_leaf_270_wb_clk_i),
    .Q(\soc.spi_video_ram_1.fifo_in_address[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11810_ (.D(_00010_),
    .CLK(clknet_leaf_60_wb_clk_i),
    .Q(\soc.spi_video_ram_1.fifo_read_request ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11811_ (.D(_00870_),
    .CLK(clknet_leaf_64_wb_clk_i),
    .Q(\soc.spi_video_ram_1.start_read ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11812_ (.D(_00871_),
    .CLK(clknet_leaf_63_wb_clk_i),
    .Q(\soc.spi_video_ram_1.initialized ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11813_ (.D(_00872_),
    .CLK(clknet_leaf_60_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.write_pointer[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11814_ (.D(_00873_),
    .CLK(clknet_leaf_48_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.write_pointer[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11815_ (.D(_00874_),
    .CLK(clknet_leaf_48_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.write_pointer[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11816_ (.D(_00875_),
    .CLK(clknet_leaf_48_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.write_pointer[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11817_ (.D(_00876_),
    .CLK(clknet_leaf_60_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.write_pointer[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11818_ (.D(_00877_),
    .CLK(clknet_leaf_61_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.read_pointer[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11819_ (.D(_00878_),
    .CLK(clknet_leaf_71_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.read_pointer[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11820_ (.D(_00879_),
    .CLK(clknet_leaf_47_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.read_pointer[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11821_ (.D(_00880_),
    .CLK(clknet_leaf_32_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.read_pointer[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11822_ (.D(_00881_),
    .CLK(clknet_leaf_32_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.read_pointer[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11823_ (.D(_00882_),
    .CLK(clknet_leaf_96_wb_clk_i),
    .Q(\soc.rom_encoder_0.input_bits_left[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11824_ (.D(_00883_),
    .CLK(clknet_leaf_96_wb_clk_i),
    .Q(\soc.rom_encoder_0.input_bits_left[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11825_ (.D(_00884_),
    .CLK(clknet_leaf_96_wb_clk_i),
    .Q(\soc.rom_encoder_0.input_bits_left[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11826_ (.D(_00885_),
    .CLK(clknet_leaf_125_wb_clk_i),
    .Q(\soc.rom_encoder_0.input_buffer[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11827_ (.D(_00886_),
    .CLK(clknet_leaf_102_wb_clk_i),
    .Q(\soc.rom_encoder_0.input_buffer[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11828_ (.D(_00887_),
    .CLK(clknet_leaf_124_wb_clk_i),
    .Q(\soc.rom_encoder_0.input_buffer[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11829_ (.D(_00888_),
    .CLK(clknet_leaf_121_wb_clk_i),
    .Q(\soc.rom_encoder_0.input_buffer[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11830_ (.D(_00889_),
    .CLK(clknet_leaf_123_wb_clk_i),
    .Q(\soc.rom_encoder_0.input_buffer[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11831_ (.D(_00890_),
    .CLK(clknet_leaf_122_wb_clk_i),
    .Q(\soc.rom_encoder_0.input_buffer[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11832_ (.D(_00891_),
    .CLK(clknet_leaf_125_wb_clk_i),
    .Q(\soc.rom_encoder_0.input_buffer[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11833_ (.D(_00892_),
    .CLK(clknet_leaf_122_wb_clk_i),
    .Q(\soc.rom_encoder_0.input_buffer[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11834_ (.D(_00893_),
    .CLK(clknet_leaf_123_wb_clk_i),
    .Q(\soc.rom_encoder_0.input_buffer[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11835_ (.D(_00894_),
    .CLK(clknet_leaf_122_wb_clk_i),
    .Q(\soc.rom_encoder_0.input_buffer[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11836_ (.D(_00895_),
    .CLK(clknet_leaf_125_wb_clk_i),
    .Q(\soc.rom_encoder_0.input_buffer[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11837_ (.D(_00896_),
    .CLK(clknet_leaf_123_wb_clk_i),
    .Q(\soc.rom_encoder_0.input_buffer[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11838_ (.D(_00897_),
    .CLK(clknet_leaf_101_wb_clk_i),
    .Q(\soc.rom_encoder_0.request_write ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11839_ (.D(_00898_),
    .CLK(clknet_leaf_102_wb_clk_i),
    .Q(\soc.rom_encoder_0.request_data_out[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11840_ (.D(_00899_),
    .CLK(clknet_5_11_0_wb_clk_i),
    .Q(\soc.rom_encoder_0.request_data_out[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11841_ (.D(_00900_),
    .CLK(clknet_leaf_170_wb_clk_i),
    .Q(\soc.rom_encoder_0.request_data_out[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11842_ (.D(_00901_),
    .CLK(clknet_leaf_170_wb_clk_i),
    .Q(\soc.rom_encoder_0.request_data_out[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11843_ (.D(_00902_),
    .CLK(clknet_leaf_95_wb_clk_i),
    .Q(\soc.rom_encoder_0.request_data_out[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11844_ (.D(_00903_),
    .CLK(clknet_leaf_95_wb_clk_i),
    .Q(\soc.rom_encoder_0.request_data_out[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11845_ (.D(_00904_),
    .CLK(clknet_leaf_169_wb_clk_i),
    .Q(\soc.rom_encoder_0.request_data_out[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11846_ (.D(_00905_),
    .CLK(clknet_leaf_166_wb_clk_i),
    .Q(\soc.rom_encoder_0.request_data_out[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11847_ (.D(_00906_),
    .CLK(clknet_leaf_169_wb_clk_i),
    .Q(\soc.rom_encoder_0.request_data_out[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11848_ (.D(_00907_),
    .CLK(clknet_leaf_122_wb_clk_i),
    .Q(\soc.rom_encoder_0.request_data_out[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11849_ (.D(_00908_),
    .CLK(clknet_leaf_87_wb_clk_i),
    .Q(\soc.rom_encoder_0.request_data_out[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11850_ (.D(_00909_),
    .CLK(clknet_leaf_107_wb_clk_i),
    .Q(\soc.rom_encoder_0.request_data_out[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11851_ (.D(_00910_),
    .CLK(clknet_leaf_93_wb_clk_i),
    .Q(\soc.rom_encoder_0.request_data_out[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11852_ (.D(_00911_),
    .CLK(clknet_leaf_106_wb_clk_i),
    .Q(\soc.rom_encoder_0.request_data_out[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11853_ (.D(_00912_),
    .CLK(clknet_leaf_100_wb_clk_i),
    .Q(\soc.rom_encoder_0.request_data_out[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11854_ (.D(_00913_),
    .CLK(clknet_leaf_96_wb_clk_i),
    .Q(\soc.rom_encoder_0.request_data_out[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11855_ (.D(_00914_),
    .CLK(clknet_leaf_92_wb_clk_i),
    .Q(\soc.rom_encoder_0.request_address[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11856_ (.D(_00915_),
    .CLK(clknet_leaf_107_wb_clk_i),
    .Q(\soc.rom_encoder_0.request_address[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11857_ (.D(_00916_),
    .CLK(clknet_leaf_92_wb_clk_i),
    .Q(\soc.rom_encoder_0.request_address[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11858_ (.D(_00917_),
    .CLK(clknet_leaf_108_wb_clk_i),
    .Q(\soc.rom_encoder_0.request_address[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11859_ (.D(_00918_),
    .CLK(clknet_leaf_106_wb_clk_i),
    .Q(\soc.rom_encoder_0.request_address[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11860_ (.D(_00919_),
    .CLK(clknet_leaf_106_wb_clk_i),
    .Q(\soc.rom_encoder_0.request_address[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11861_ (.D(_00920_),
    .CLK(clknet_leaf_105_wb_clk_i),
    .Q(\soc.rom_encoder_0.request_address[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11862_ (.D(_00921_),
    .CLK(clknet_leaf_109_wb_clk_i),
    .Q(\soc.rom_encoder_0.request_address[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11863_ (.D(_00922_),
    .CLK(clknet_leaf_105_wb_clk_i),
    .Q(\soc.rom_encoder_0.request_address[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11864_ (.D(_00923_),
    .CLK(clknet_leaf_109_wb_clk_i),
    .Q(\soc.rom_encoder_0.request_address[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11865_ (.D(_00924_),
    .CLK(clknet_leaf_109_wb_clk_i),
    .Q(\soc.rom_encoder_0.request_address[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11866_ (.D(_00925_),
    .CLK(clknet_leaf_104_wb_clk_i),
    .Q(\soc.rom_encoder_0.request_address[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11867_ (.D(_00926_),
    .CLK(clknet_leaf_104_wb_clk_i),
    .Q(\soc.rom_encoder_0.request_address[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11868_ (.D(_00927_),
    .CLK(clknet_5_15_0_wb_clk_i),
    .Q(\soc.rom_encoder_0.request_address[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11869_ (.D(_00928_),
    .CLK(clknet_leaf_102_wb_clk_i),
    .Q(\soc.rom_encoder_0.request_address[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11870_ (.D(_00929_),
    .CLK(clknet_leaf_165_wb_clk_i),
    .Q(net58));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11871_ (.D(_00930_),
    .CLK(clknet_leaf_165_wb_clk_i),
    .Q(net59));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11872_ (.D(_00931_),
    .CLK(clknet_leaf_165_wb_clk_i),
    .Q(net60));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11873_ (.D(_00932_),
    .CLK(clknet_leaf_165_wb_clk_i),
    .Q(net61));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11874_ (.D(_00933_),
    .CLK(clknet_leaf_221_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[3][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11875_ (.D(_00934_),
    .CLK(clknet_leaf_215_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[3][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11876_ (.D(_00935_),
    .CLK(clknet_leaf_258_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[3][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11877_ (.D(_00936_),
    .CLK(clknet_leaf_259_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[3][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11878_ (.D(_00937_),
    .CLK(clknet_leaf_199_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[3][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11879_ (.D(_00938_),
    .CLK(clknet_leaf_214_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[3][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11880_ (.D(_00939_),
    .CLK(clknet_leaf_247_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[3][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11881_ (.D(_00940_),
    .CLK(clknet_5_19_0_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[3][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11882_ (.D(_00941_),
    .CLK(clknet_leaf_216_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[3][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11883_ (.D(_00942_),
    .CLK(clknet_leaf_249_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[3][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11884_ (.D(_00943_),
    .CLK(clknet_leaf_17_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[3][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11885_ (.D(_00944_),
    .CLK(clknet_leaf_14_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[3][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11886_ (.D(_00945_),
    .CLK(clknet_leaf_1_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[3][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11887_ (.D(_00946_),
    .CLK(clknet_leaf_320_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[3][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11888_ (.D(_00947_),
    .CLK(clknet_leaf_318_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[3][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11889_ (.D(_00948_),
    .CLK(clknet_leaf_320_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[3][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11890_ (.D(_00949_),
    .CLK(clknet_leaf_25_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[3][16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11891_ (.D(_00950_),
    .CLK(clknet_leaf_78_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[3][17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11892_ (.D(_00951_),
    .CLK(clknet_leaf_77_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[3][18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11893_ (.D(_00952_),
    .CLK(clknet_leaf_74_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[3][19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11894_ (.D(_00953_),
    .CLK(clknet_leaf_45_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[3][20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11895_ (.D(_00954_),
    .CLK(clknet_leaf_230_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[3][21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11896_ (.D(_00955_),
    .CLK(clknet_leaf_253_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[3][22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11897_ (.D(_00956_),
    .CLK(clknet_leaf_241_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[3][23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11898_ (.D(_00957_),
    .CLK(clknet_leaf_298_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[3][24] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11899_ (.D(_00958_),
    .CLK(clknet_leaf_234_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[3][25] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11900_ (.D(_00959_),
    .CLK(clknet_leaf_296_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[3][26] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11901_ (.D(_00960_),
    .CLK(clknet_leaf_44_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[3][27] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11902_ (.D(_00961_),
    .CLK(clknet_leaf_296_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[3][28] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11903_ (.D(_00962_),
    .CLK(clknet_leaf_99_wb_clk_i),
    .Q(\soc.rom_encoder_0.initialized ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11904_ (.D(_00963_),
    .CLK(clknet_leaf_124_wb_clk_i),
    .Q(\soc.cpu.DMuxJMP.sel[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11905_ (.D(_00964_),
    .CLK(clknet_leaf_127_wb_clk_i),
    .Q(\soc.cpu.DMuxJMP.sel[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11906_ (.D(_00965_),
    .CLK(clknet_leaf_124_wb_clk_i),
    .Q(\soc.cpu.DMuxJMP.sel[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11907_ (.D(_00966_),
    .CLK(clknet_leaf_121_wb_clk_i),
    .Q(\soc.cpu.instruction[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11908_ (.D(_00967_),
    .CLK(clknet_leaf_127_wb_clk_i),
    .Q(\soc.cpu.instruction[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11909_ (.D(_00968_),
    .CLK(clknet_leaf_121_wb_clk_i),
    .Q(\soc.cpu.instruction[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11910_ (.D(_00969_),
    .CLK(clknet_leaf_128_wb_clk_i),
    .Q(\soc.cpu.ALU.no ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11911_ (.D(_00970_),
    .CLK(clknet_leaf_127_wb_clk_i),
    .Q(\soc.cpu.ALU.f ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11912_ (.D(_00971_),
    .CLK(clknet_5_13_0_wb_clk_i),
    .Q(\soc.cpu.ALU.ny ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11913_ (.D(_00972_),
    .CLK(clknet_5_26_0_wb_clk_i),
    .Q(\soc.cpu.ALU.zy ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11914_ (.D(_00973_),
    .CLK(clknet_leaf_128_wb_clk_i),
    .Q(\soc.cpu.ALU.nx ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11915_ (.D(_00974_),
    .CLK(clknet_leaf_121_wb_clk_i),
    .Q(\soc.cpu.ALU.zx ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11916_ (.D(_00975_),
    .CLK(clknet_leaf_119_wb_clk_i),
    .Q(\soc.cpu.instruction[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11917_ (.D(_00976_),
    .CLK(clknet_leaf_122_wb_clk_i),
    .Q(\soc.cpu.instruction[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11918_ (.D(_00977_),
    .CLK(clknet_leaf_121_wb_clk_i),
    .Q(\soc.cpu.instruction[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11919_ (.D(_00978_),
    .CLK(clknet_leaf_121_wb_clk_i),
    .Q(\soc.cpu.instruction[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11920_ (.D(_00979_),
    .CLK(clknet_leaf_99_wb_clk_i),
    .Q(net62));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11921_ (.D(_00980_),
    .CLK(clknet_leaf_100_wb_clk_i),
    .Q(\soc.rom_encoder_0.sram_sio_oe ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11922_ (.D(_00981_),
    .CLK(clknet_leaf_97_wb_clk_i),
    .Q(\soc.rom_encoder_0.current_state[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11923_ (.D(_00982_),
    .CLK(clknet_leaf_97_wb_clk_i),
    .Q(\soc.rom_encoder_0.current_state[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11924_ (.D(_00983_),
    .CLK(clknet_leaf_98_wb_clk_i),
    .Q(\soc.rom_encoder_0.current_state[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11925_ (.D(_00984_),
    .CLK(clknet_leaf_86_wb_clk_i),
    .Q(\soc.rom_encoder_0.initializing_step[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11926_ (.D(_00985_),
    .CLK(clknet_leaf_97_wb_clk_i),
    .Q(\soc.rom_encoder_0.initializing_step[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11927_ (.D(_00986_),
    .CLK(clknet_leaf_86_wb_clk_i),
    .Q(\soc.rom_encoder_0.initializing_step[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11928_ (.D(_00987_),
    .CLK(clknet_leaf_85_wb_clk_i),
    .Q(\soc.rom_encoder_0.initializing_step[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11929_ (.D(_00988_),
    .CLK(clknet_leaf_86_wb_clk_i),
    .Q(\soc.rom_encoder_0.initializing_step[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11930_ (.D(_00989_),
    .CLK(clknet_leaf_160_wb_clk_i),
    .Q(\soc.ram_encoder_0.toggled_sram_sck ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11931_ (.D(_00990_),
    .CLK(clknet_leaf_164_wb_clk_i),
    .Q(\soc.ram_encoder_0.input_bits_left[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11932_ (.D(_00991_),
    .CLK(clknet_leaf_164_wb_clk_i),
    .Q(\soc.ram_encoder_0.input_bits_left[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11933_ (.D(_00992_),
    .CLK(clknet_leaf_165_wb_clk_i),
    .Q(\soc.ram_encoder_0.input_bits_left[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11934_ (.D(_00993_),
    .CLK(clknet_leaf_158_wb_clk_i),
    .Q(\soc.ram_encoder_0.input_buffer[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11935_ (.D(_00994_),
    .CLK(clknet_leaf_158_wb_clk_i),
    .Q(\soc.ram_encoder_0.input_buffer[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11936_ (.D(_00995_),
    .CLK(clknet_leaf_160_wb_clk_i),
    .Q(\soc.ram_encoder_0.input_buffer[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11937_ (.D(_00996_),
    .CLK(clknet_leaf_157_wb_clk_i),
    .Q(\soc.ram_encoder_0.input_buffer[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11938_ (.D(_00997_),
    .CLK(clknet_leaf_158_wb_clk_i),
    .Q(\soc.ram_encoder_0.input_buffer[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11939_ (.D(_00998_),
    .CLK(clknet_leaf_158_wb_clk_i),
    .Q(\soc.ram_encoder_0.input_buffer[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11940_ (.D(_00999_),
    .CLK(clknet_leaf_160_wb_clk_i),
    .Q(\soc.ram_encoder_0.input_buffer[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11941_ (.D(_01000_),
    .CLK(clknet_leaf_159_wb_clk_i),
    .Q(\soc.ram_encoder_0.input_buffer[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11942_ (.D(_01001_),
    .CLK(clknet_leaf_159_wb_clk_i),
    .Q(\soc.ram_encoder_0.input_buffer[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11943_ (.D(_01002_),
    .CLK(clknet_leaf_159_wb_clk_i),
    .Q(\soc.ram_encoder_0.input_buffer[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11944_ (.D(_01003_),
    .CLK(clknet_leaf_160_wb_clk_i),
    .Q(\soc.ram_encoder_0.input_buffer[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11945_ (.D(_01004_),
    .CLK(clknet_leaf_161_wb_clk_i),
    .Q(\soc.ram_encoder_0.input_buffer[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11946_ (.D(_01005_),
    .CLK(clknet_leaf_154_wb_clk_i),
    .Q(\soc.ram_encoder_0.request_write ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11947_ (.D(_01006_),
    .CLK(clknet_leaf_152_wb_clk_i),
    .Q(\soc.ram_encoder_0.request_data_out[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11948_ (.D(_01007_),
    .CLK(clknet_leaf_148_wb_clk_i),
    .Q(\soc.ram_encoder_0.request_data_out[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11949_ (.D(_01008_),
    .CLK(clknet_leaf_156_wb_clk_i),
    .Q(\soc.ram_encoder_0.request_data_out[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11950_ (.D(_01009_),
    .CLK(clknet_leaf_156_wb_clk_i),
    .Q(\soc.ram_encoder_0.request_data_out[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11951_ (.D(_01010_),
    .CLK(clknet_leaf_155_wb_clk_i),
    .Q(\soc.ram_encoder_0.request_data_out[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11952_ (.D(_01011_),
    .CLK(clknet_leaf_153_wb_clk_i),
    .Q(\soc.ram_encoder_0.request_data_out[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11953_ (.D(_01012_),
    .CLK(clknet_leaf_152_wb_clk_i),
    .Q(\soc.ram_encoder_0.request_data_out[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11954_ (.D(_01013_),
    .CLK(clknet_leaf_153_wb_clk_i),
    .Q(\soc.ram_encoder_0.request_data_out[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11955_ (.D(_01014_),
    .CLK(clknet_leaf_154_wb_clk_i),
    .Q(\soc.ram_encoder_0.request_data_out[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11956_ (.D(_01015_),
    .CLK(clknet_leaf_154_wb_clk_i),
    .Q(\soc.ram_encoder_0.request_data_out[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11957_ (.D(_01016_),
    .CLK(clknet_leaf_159_wb_clk_i),
    .Q(\soc.ram_encoder_0.request_data_out[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11958_ (.D(_01017_),
    .CLK(clknet_leaf_118_wb_clk_i),
    .Q(\soc.ram_encoder_0.request_data_out[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11959_ (.D(_01018_),
    .CLK(clknet_leaf_114_wb_clk_i),
    .Q(\soc.ram_encoder_0.request_data_out[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11960_ (.D(_01019_),
    .CLK(clknet_leaf_162_wb_clk_i),
    .Q(\soc.ram_encoder_0.request_data_out[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11961_ (.D(_01020_),
    .CLK(clknet_leaf_114_wb_clk_i),
    .Q(\soc.ram_encoder_0.request_data_out[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11962_ (.D(_01021_),
    .CLK(clknet_leaf_162_wb_clk_i),
    .Q(\soc.ram_encoder_0.request_data_out[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11963_ (.D(_01022_),
    .CLK(clknet_leaf_148_wb_clk_i),
    .Q(\soc.ram_encoder_0.request_address[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11964_ (.D(_01023_),
    .CLK(clknet_leaf_149_wb_clk_i),
    .Q(\soc.ram_encoder_0.request_address[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11965_ (.D(_01024_),
    .CLK(clknet_leaf_147_wb_clk_i),
    .Q(\soc.ram_encoder_0.request_address[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11966_ (.D(_01025_),
    .CLK(clknet_leaf_146_wb_clk_i),
    .Q(\soc.ram_encoder_0.request_address[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11967_ (.D(_01026_),
    .CLK(clknet_leaf_147_wb_clk_i),
    .Q(\soc.ram_encoder_0.request_address[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11968_ (.D(_01027_),
    .CLK(clknet_leaf_183_wb_clk_i),
    .Q(\soc.ram_encoder_0.request_address[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11969_ (.D(_01028_),
    .CLK(clknet_leaf_183_wb_clk_i),
    .Q(\soc.ram_encoder_0.request_address[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11970_ (.D(_01029_),
    .CLK(clknet_leaf_147_wb_clk_i),
    .Q(\soc.ram_encoder_0.request_address[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11971_ (.D(_01030_),
    .CLK(clknet_leaf_148_wb_clk_i),
    .Q(\soc.ram_encoder_0.request_address[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11972_ (.D(_01031_),
    .CLK(clknet_leaf_150_wb_clk_i),
    .Q(\soc.ram_encoder_0.request_address[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11973_ (.D(_01032_),
    .CLK(clknet_leaf_169_wb_clk_i),
    .Q(\soc.ram_encoder_0.request_address[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11974_ (.D(_01033_),
    .CLK(clknet_leaf_153_wb_clk_i),
    .Q(\soc.ram_encoder_0.request_address[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11975_ (.D(_01034_),
    .CLK(clknet_leaf_168_wb_clk_i),
    .Q(\soc.ram_encoder_0.request_address[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11976_ (.D(_01035_),
    .CLK(clknet_leaf_153_wb_clk_i),
    .Q(\soc.ram_encoder_0.request_address[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11977_ (.D(_01036_),
    .CLK(clknet_leaf_153_wb_clk_i),
    .Q(\soc.ram_encoder_0.request_address[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11978_ (.D(_01037_),
    .CLK(clknet_leaf_127_wb_clk_i),
    .Q(\soc.ram_encoder_0.initialized ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11979_ (.D(_01038_),
    .CLK(clknet_leaf_157_wb_clk_i),
    .Q(\soc.ram_data_out[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11980_ (.D(_01039_),
    .CLK(clknet_leaf_157_wb_clk_i),
    .Q(\soc.ram_data_out[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11981_ (.D(_01040_),
    .CLK(clknet_leaf_156_wb_clk_i),
    .Q(\soc.ram_data_out[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11982_ (.D(_01041_),
    .CLK(clknet_leaf_157_wb_clk_i),
    .Q(\soc.ram_data_out[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11983_ (.D(_01042_),
    .CLK(clknet_leaf_158_wb_clk_i),
    .Q(\soc.ram_data_out[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11984_ (.D(_01043_),
    .CLK(clknet_leaf_155_wb_clk_i),
    .Q(\soc.ram_data_out[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11985_ (.D(_01044_),
    .CLK(clknet_leaf_144_wb_clk_i),
    .Q(\soc.ram_data_out[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11986_ (.D(_01045_),
    .CLK(clknet_leaf_144_wb_clk_i),
    .Q(\soc.ram_data_out[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11987_ (.D(_01046_),
    .CLK(clknet_leaf_158_wb_clk_i),
    .Q(\soc.ram_data_out[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11988_ (.D(_01047_),
    .CLK(clknet_leaf_158_wb_clk_i),
    .Q(\soc.ram_data_out[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11989_ (.D(_01048_),
    .CLK(clknet_leaf_118_wb_clk_i),
    .Q(\soc.ram_data_out[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11990_ (.D(_01049_),
    .CLK(clknet_leaf_119_wb_clk_i),
    .Q(\soc.ram_data_out[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11991_ (.D(_01050_),
    .CLK(clknet_leaf_118_wb_clk_i),
    .Q(\soc.ram_data_out[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11992_ (.D(_01051_),
    .CLK(clknet_leaf_118_wb_clk_i),
    .Q(\soc.ram_data_out[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11993_ (.D(_01052_),
    .CLK(clknet_leaf_117_wb_clk_i),
    .Q(\soc.ram_data_out[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11994_ (.D(_01053_),
    .CLK(clknet_leaf_118_wb_clk_i),
    .Q(\soc.ram_data_out[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11995_ (.D(_01054_),
    .CLK(clknet_leaf_161_wb_clk_i),
    .Q(net81));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11996_ (.D(_01055_),
    .CLK(clknet_leaf_161_wb_clk_i),
    .Q(\soc.ram_encoder_0.sram_sio_oe ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11997_ (.D(_01056_),
    .CLK(clknet_leaf_161_wb_clk_i),
    .Q(\soc.ram_encoder_0.current_state[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11998_ (.D(_01057_),
    .CLK(clknet_leaf_165_wb_clk_i),
    .Q(\soc.ram_encoder_0.current_state[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11999_ (.D(_01058_),
    .CLK(clknet_leaf_164_wb_clk_i),
    .Q(\soc.ram_encoder_0.current_state[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12000_ (.D(_01059_),
    .CLK(clknet_leaf_163_wb_clk_i),
    .Q(\soc.ram_encoder_0.initializing_step[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12001_ (.D(_01060_),
    .CLK(clknet_leaf_163_wb_clk_i),
    .Q(\soc.ram_encoder_0.initializing_step[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12002_ (.D(_01061_),
    .CLK(clknet_leaf_163_wb_clk_i),
    .Q(\soc.ram_encoder_0.initializing_step[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12003_ (.D(_01062_),
    .CLK(clknet_leaf_163_wb_clk_i),
    .Q(\soc.ram_encoder_0.initializing_step[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12004_ (.D(_01063_),
    .CLK(clknet_leaf_164_wb_clk_i),
    .Q(\soc.ram_encoder_0.initializing_step[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12005_ (.D(_01064_),
    .CLK(clknet_leaf_115_wb_clk_i),
    .Q(\soc.hack_clock_0.counter[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12006_ (.D(_01065_),
    .CLK(clknet_leaf_113_wb_clk_i),
    .Q(\soc.hack_clock_0.counter[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12007_ (.D(_01066_),
    .CLK(clknet_leaf_113_wb_clk_i),
    .Q(\soc.hack_clock_0.counter[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12008_ (.D(_01067_),
    .CLK(clknet_leaf_163_wb_clk_i),
    .Q(\soc.hack_clock_0.counter[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12009_ (.D(_01068_),
    .CLK(clknet_leaf_163_wb_clk_i),
    .Q(\soc.hack_clock_0.counter[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12010_ (.D(_01069_),
    .CLK(clknet_leaf_113_wb_clk_i),
    .Q(\soc.hack_clock_0.counter[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12011_ (.D(_01070_),
    .CLK(clknet_leaf_113_wb_clk_i),
    .Q(\soc.hack_clock_0.counter[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12012_ (.D(_01071_),
    .CLK(clknet_leaf_212_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[5][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12013_ (.D(_01072_),
    .CLK(clknet_leaf_214_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[5][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12014_ (.D(_01073_),
    .CLK(clknet_leaf_266_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[5][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12015_ (.D(_01074_),
    .CLK(clknet_leaf_265_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[5][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12016_ (.D(_01075_),
    .CLK(clknet_leaf_254_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[5][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12017_ (.D(_01076_),
    .CLK(clknet_leaf_227_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[5][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12018_ (.D(_01077_),
    .CLK(clknet_leaf_246_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[5][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12019_ (.D(_01078_),
    .CLK(clknet_leaf_243_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[5][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12020_ (.D(_01079_),
    .CLK(clknet_leaf_228_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[5][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12021_ (.D(_01080_),
    .CLK(clknet_leaf_246_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[5][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12022_ (.D(_01081_),
    .CLK(clknet_leaf_15_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[5][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12023_ (.D(_01082_),
    .CLK(clknet_leaf_38_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[5][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12024_ (.D(_01083_),
    .CLK(clknet_leaf_309_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[5][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12025_ (.D(_01084_),
    .CLK(clknet_leaf_312_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[5][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12026_ (.D(_01085_),
    .CLK(clknet_leaf_313_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[5][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12027_ (.D(_01086_),
    .CLK(clknet_leaf_312_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[5][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12028_ (.D(_01087_),
    .CLK(clknet_leaf_74_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[5][16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12029_ (.D(_01088_),
    .CLK(clknet_leaf_67_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[5][17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12030_ (.D(_01089_),
    .CLK(clknet_leaf_67_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[5][18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12031_ (.D(_01090_),
    .CLK(clknet_leaf_72_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[5][19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12032_ (.D(_01091_),
    .CLK(clknet_leaf_59_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[5][20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12033_ (.D(_01092_),
    .CLK(clknet_leaf_292_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[5][21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12034_ (.D(_01093_),
    .CLK(clknet_leaf_270_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[5][22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12035_ (.D(_01094_),
    .CLK(clknet_leaf_287_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[5][23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12036_ (.D(_01095_),
    .CLK(clknet_leaf_302_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[5][24] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12037_ (.D(_01096_),
    .CLK(clknet_leaf_289_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[5][25] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12038_ (.D(_01097_),
    .CLK(clknet_leaf_295_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[5][26] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12039_ (.D(_01098_),
    .CLK(clknet_leaf_273_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[5][27] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12040_ (.D(_01099_),
    .CLK(clknet_leaf_274_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[5][28] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12041_ (.D(_01100_),
    .CLK(clknet_leaf_99_wb_clk_i),
    .Q(\soc.rom_loader.rom_request ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12042_ (.D(_01101_),
    .CLK(clknet_leaf_125_wb_clk_i),
    .Q(\soc.rom_loader.writing ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12043_ (.D(net20),
    .CLK(clknet_leaf_297_wb_clk_i),
    .Q(\soc.rom_encoder_0.data_out[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12044_ (.D(net21),
    .CLK(clknet_leaf_87_wb_clk_i),
    .Q(\soc.rom_encoder_0.data_out[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12045_ (.D(net22),
    .CLK(clknet_5_31_0_wb_clk_i),
    .Q(\soc.rom_encoder_0.data_out[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12046_ (.D(net23),
    .CLK(clknet_5_31_0_wb_clk_i),
    .Q(\soc.rom_encoder_0.data_out[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12047_ (.D(net24),
    .CLK(clknet_leaf_95_wb_clk_i),
    .Q(\soc.rom_encoder_0.data_out[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12048_ (.D(net25),
    .CLK(clknet_opt_1_0_wb_clk_i),
    .Q(\soc.rom_encoder_0.data_out[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12049_ (.D(net26),
    .CLK(clknet_leaf_173_wb_clk_i),
    .Q(\soc.rom_encoder_0.data_out[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12050_ (.D(net27),
    .CLK(clknet_5_31_0_wb_clk_i),
    .Q(\soc.rom_encoder_0.data_out[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12051_ (.D(net28),
    .CLK(clknet_5_31_0_wb_clk_i),
    .Q(\soc.rom_encoder_0.data_out[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12052_ (.D(net30),
    .CLK(clknet_leaf_112_wb_clk_i),
    .Q(\soc.rom_encoder_0.data_out[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12053_ (.D(net31),
    .CLK(clknet_leaf_87_wb_clk_i),
    .Q(\soc.rom_encoder_0.data_out[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12054_ (.D(net32),
    .CLK(clknet_leaf_108_wb_clk_i),
    .Q(\soc.rom_encoder_0.data_out[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12055_ (.D(net33),
    .CLK(clknet_opt_2_0_wb_clk_i),
    .Q(\soc.rom_encoder_0.data_out[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12056_ (.D(net34),
    .CLK(clknet_leaf_106_wb_clk_i),
    .Q(\soc.rom_encoder_0.data_out[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12057_ (.D(net35),
    .CLK(clknet_leaf_173_wb_clk_i),
    .Q(\soc.rom_encoder_0.data_out[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12058_ (.D(net36),
    .CLK(clknet_leaf_315_wb_clk_i),
    .Q(\soc.rom_encoder_0.data_out[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _12059_ (.D(_01102_),
    .CLK(clknet_leaf_99_wb_clk_i),
    .Q(\soc.rom_encoder_0.toggled_sram_sck ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12060_ (.D(_01103_),
    .CLK(clknet_leaf_107_wb_clk_i),
    .Q(\soc.rom_loader.current_address[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12061_ (.D(_01104_),
    .CLK(clknet_leaf_107_wb_clk_i),
    .Q(\soc.rom_loader.current_address[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12062_ (.D(_01105_),
    .CLK(clknet_leaf_108_wb_clk_i),
    .Q(\soc.rom_loader.current_address[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12063_ (.D(_01106_),
    .CLK(clknet_leaf_112_wb_clk_i),
    .Q(\soc.rom_loader.current_address[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12064_ (.D(_01107_),
    .CLK(clknet_leaf_112_wb_clk_i),
    .Q(\soc.rom_loader.current_address[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12065_ (.D(_01108_),
    .CLK(clknet_leaf_112_wb_clk_i),
    .Q(\soc.rom_loader.current_address[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12066_ (.D(_01109_),
    .CLK(clknet_leaf_108_wb_clk_i),
    .Q(\soc.rom_loader.current_address[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12067_ (.D(_01110_),
    .CLK(clknet_leaf_111_wb_clk_i),
    .Q(\soc.rom_loader.current_address[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12068_ (.D(_01111_),
    .CLK(clknet_leaf_111_wb_clk_i),
    .Q(\soc.rom_loader.current_address[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12069_ (.D(_01112_),
    .CLK(clknet_leaf_111_wb_clk_i),
    .Q(\soc.rom_loader.current_address[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12070_ (.D(_01113_),
    .CLK(clknet_leaf_109_wb_clk_i),
    .Q(\soc.rom_loader.current_address[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12071_ (.D(_01114_),
    .CLK(clknet_leaf_110_wb_clk_i),
    .Q(\soc.rom_loader.current_address[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12072_ (.D(_01115_),
    .CLK(clknet_leaf_109_wb_clk_i),
    .Q(\soc.rom_loader.current_address[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12073_ (.D(_01116_),
    .CLK(clknet_leaf_102_wb_clk_i),
    .Q(\soc.rom_loader.current_address[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12074_ (.D(_01117_),
    .CLK(clknet_leaf_110_wb_clk_i),
    .Q(\soc.rom_loader.current_address[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12075_ (.D(_01118_),
    .CLK(clknet_leaf_99_wb_clk_i),
    .Q(\soc.rom_loader.wait_fall_clk ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12076_ (.D(_01119_),
    .CLK(clknet_leaf_129_wb_clk_i),
    .Q(net83));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _12077_ (.D(\soc.cpu.PC.in[0] ),
    .CLK(net84),
    .Q(\soc.cpu.AReg.data[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _12078_ (.D(\soc.cpu.PC.in[1] ),
    .CLK(net85),
    .Q(\soc.cpu.AReg.data[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12079_ (.D(\soc.cpu.PC.in[2] ),
    .CLK(net84),
    .Q(\soc.cpu.AReg.data[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12080_ (.D(\soc.cpu.PC.in[3] ),
    .CLK(net84),
    .Q(\soc.cpu.AReg.data[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12081_ (.D(\soc.cpu.PC.in[4] ),
    .CLK(net84),
    .Q(\soc.cpu.AReg.data[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _12082_ (.D(\soc.cpu.PC.in[5] ),
    .CLK(net89),
    .Q(\soc.cpu.AReg.data[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12083_ (.D(\soc.cpu.PC.in[6] ),
    .CLK(net84),
    .Q(\soc.cpu.AReg.data[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12084_ (.D(\soc.cpu.PC.in[7] ),
    .CLK(net84),
    .Q(\soc.cpu.AReg.data[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12085_ (.D(\soc.cpu.PC.in[8] ),
    .CLK(net84),
    .Q(\soc.cpu.AReg.data[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12086_ (.D(\soc.cpu.PC.in[9] ),
    .CLK(net90),
    .Q(\soc.cpu.AReg.data[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _12087_ (.D(\soc.cpu.PC.in[10] ),
    .CLK(net84),
    .Q(\soc.cpu.AReg.data[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _12088_ (.D(\soc.cpu.PC.in[11] ),
    .CLK(net84),
    .Q(\soc.cpu.AReg.data[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _12089_ (.D(\soc.cpu.PC.in[12] ),
    .CLK(net89),
    .Q(\soc.cpu.AReg.data[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _12090_ (.D(\soc.cpu.PC.in[13] ),
    .CLK(net89),
    .Q(\soc.cpu.AReg.data[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _12091_ (.D(\soc.cpu.PC.in[14] ),
    .CLK(net89),
    .Q(\soc.cpu.AReg.data[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12092_ (.D(_01120_),
    .CLK(net86),
    .Q(\soc.cpu.ALU.x[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12093_ (.D(_01121_),
    .CLK(net86),
    .Q(\soc.cpu.ALU.x[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12094_ (.D(_01122_),
    .CLK(net86),
    .Q(\soc.cpu.ALU.x[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12095_ (.D(_01123_),
    .CLK(net86),
    .Q(\soc.cpu.ALU.x[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12096_ (.D(_01124_),
    .CLK(net86),
    .Q(\soc.cpu.ALU.x[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12097_ (.D(_01125_),
    .CLK(net86),
    .Q(\soc.cpu.ALU.x[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12098_ (.D(_01126_),
    .CLK(net86),
    .Q(\soc.cpu.ALU.x[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12099_ (.D(_01127_),
    .CLK(net86),
    .Q(\soc.cpu.ALU.x[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12100_ (.D(_01128_),
    .CLK(net85),
    .Q(\soc.cpu.ALU.x[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12101_ (.D(_01129_),
    .CLK(net85),
    .Q(\soc.cpu.ALU.x[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12102_ (.D(_01130_),
    .CLK(net85),
    .Q(\soc.cpu.ALU.x[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12103_ (.D(_01131_),
    .CLK(net85),
    .Q(\soc.cpu.ALU.x[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12104_ (.D(_01132_),
    .CLK(net85),
    .Q(\soc.cpu.ALU.x[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12105_ (.D(_01133_),
    .CLK(net85),
    .Q(\soc.cpu.ALU.x[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12106_ (.D(_01134_),
    .CLK(net85),
    .Q(\soc.cpu.ALU.x[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12107_ (.D(_01135_),
    .CLK(net85),
    .Q(\soc.cpu.ALU.x[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12108_ (.D(_01136_),
    .CLK(clknet_leaf_245_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[6][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12109_ (.D(_01137_),
    .CLK(clknet_leaf_245_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[6][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12110_ (.D(_01138_),
    .CLK(clknet_leaf_265_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[6][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12111_ (.D(_01139_),
    .CLK(clknet_leaf_266_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[6][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12112_ (.D(_01140_),
    .CLK(clknet_leaf_266_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[6][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12113_ (.D(_01141_),
    .CLK(clknet_leaf_245_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[6][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12114_ (.D(_01142_),
    .CLK(clknet_leaf_246_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[6][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12115_ (.D(_01143_),
    .CLK(clknet_leaf_243_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[6][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12116_ (.D(_01144_),
    .CLK(clknet_leaf_244_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[6][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12117_ (.D(_01145_),
    .CLK(clknet_leaf_249_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[6][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12118_ (.D(_01146_),
    .CLK(clknet_leaf_15_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[6][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12119_ (.D(_01147_),
    .CLK(clknet_leaf_40_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[6][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12120_ (.D(_01148_),
    .CLK(clknet_leaf_309_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[6][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12121_ (.D(_01149_),
    .CLK(clknet_leaf_314_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[6][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12122_ (.D(_01150_),
    .CLK(clknet_leaf_317_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[6][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12123_ (.D(_01151_),
    .CLK(clknet_leaf_316_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[6][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12124_ (.D(_01152_),
    .CLK(clknet_leaf_75_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[6][16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12125_ (.D(_01153_),
    .CLK(clknet_leaf_80_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[6][17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12126_ (.D(_01154_),
    .CLK(clknet_leaf_79_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[6][18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12127_ (.D(_01155_),
    .CLK(clknet_leaf_74_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[6][19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12128_ (.D(_01156_),
    .CLK(clknet_leaf_48_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[6][20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12129_ (.D(_01157_),
    .CLK(clknet_leaf_289_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[6][21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12130_ (.D(_01158_),
    .CLK(clknet_leaf_269_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[6][22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12131_ (.D(_01159_),
    .CLK(clknet_leaf_285_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[6][23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12132_ (.D(_01160_),
    .CLK(clknet_leaf_301_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[6][24] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12133_ (.D(_01161_),
    .CLK(clknet_leaf_289_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[6][25] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12134_ (.D(_01162_),
    .CLK(clknet_leaf_295_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[6][26] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12135_ (.D(_01163_),
    .CLK(clknet_leaf_273_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[6][27] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12136_ (.D(_01164_),
    .CLK(clknet_leaf_274_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[6][28] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12137_ (.D(_01165_),
    .CLK(clknet_leaf_163_wb_clk_i),
    .Q(\soc.cpu.AReg.clk ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12138_ (.D(_01166_),
    .CLK(net88),
    .Q(\soc.cpu.PC.REG.data[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12139_ (.D(_01167_),
    .CLK(net89),
    .Q(\soc.cpu.PC.REG.data[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12140_ (.D(_01168_),
    .CLK(net88),
    .Q(\soc.cpu.PC.REG.data[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12141_ (.D(_01169_),
    .CLK(net88),
    .Q(\soc.cpu.PC.REG.data[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12142_ (.D(_01170_),
    .CLK(net88),
    .Q(\soc.cpu.PC.REG.data[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12143_ (.D(_01171_),
    .CLK(net88),
    .Q(\soc.cpu.PC.REG.data[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12144_ (.D(_01172_),
    .CLK(net88),
    .Q(\soc.cpu.PC.REG.data[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12145_ (.D(_01173_),
    .CLK(net88),
    .Q(\soc.cpu.PC.REG.data[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12146_ (.D(_01174_),
    .CLK(net89),
    .Q(\soc.cpu.PC.REG.data[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12147_ (.D(_01175_),
    .CLK(net88),
    .Q(\soc.cpu.PC.REG.data[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12148_ (.D(_01176_),
    .CLK(net88),
    .Q(\soc.cpu.PC.REG.data[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12149_ (.D(_01177_),
    .CLK(net88),
    .Q(\soc.cpu.PC.REG.data[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12150_ (.D(_01178_),
    .CLK(net89),
    .Q(\soc.cpu.PC.REG.data[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12151_ (.D(_01179_),
    .CLK(net89),
    .Q(\soc.cpu.PC.REG.data[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12152_ (.D(_01180_),
    .CLK(net89),
    .Q(\soc.cpu.PC.REG.data[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12153_ (.D(_01181_),
    .CLK(clknet_leaf_162_wb_clk_i),
    .Q(\soc.hack_clk_strobe ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12154_ (.D(_01182_),
    .CLK(clknet_leaf_160_wb_clk_i),
    .Q(\soc.synch_hack_writeM ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12155_ (.D(_01183_),
    .CLK(clknet_leaf_144_wb_clk_i),
    .Q(\soc.ram_encoder_0.address[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12156_ (.D(_01184_),
    .CLK(clknet_leaf_144_wb_clk_i),
    .Q(\soc.ram_encoder_0.address[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12157_ (.D(_01185_),
    .CLK(clknet_leaf_147_wb_clk_i),
    .Q(\soc.ram_encoder_0.address[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12158_ (.D(_01186_),
    .CLK(clknet_leaf_145_wb_clk_i),
    .Q(\soc.ram_encoder_0.address[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12159_ (.D(_01187_),
    .CLK(clknet_leaf_145_wb_clk_i),
    .Q(\soc.ram_encoder_0.address[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12160_ (.D(_01188_),
    .CLK(clknet_leaf_149_wb_clk_i),
    .Q(\soc.ram_encoder_0.address[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12161_ (.D(_01189_),
    .CLK(clknet_leaf_185_wb_clk_i),
    .Q(\soc.ram_encoder_0.address[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12162_ (.D(_01190_),
    .CLK(clknet_leaf_146_wb_clk_i),
    .Q(\soc.ram_encoder_0.address[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12163_ (.D(_01191_),
    .CLK(clknet_leaf_148_wb_clk_i),
    .Q(\soc.ram_encoder_0.address[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12164_ (.D(_01192_),
    .CLK(clknet_leaf_151_wb_clk_i),
    .Q(\soc.ram_encoder_0.address[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12165_ (.D(_01193_),
    .CLK(clknet_leaf_151_wb_clk_i),
    .Q(\soc.ram_encoder_0.address[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12166_ (.D(_01194_),
    .CLK(clknet_leaf_153_wb_clk_i),
    .Q(\soc.ram_encoder_0.address[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12167_ (.D(_01195_),
    .CLK(clknet_leaf_168_wb_clk_i),
    .Q(\soc.ram_encoder_0.address[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12168_ (.D(_01196_),
    .CLK(clknet_leaf_152_wb_clk_i),
    .Q(\soc.ram_encoder_0.address[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12169_ (.D(_01197_),
    .CLK(clknet_leaf_154_wb_clk_i),
    .Q(\soc.ram_encoder_0.address[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12170_ (.D(_01198_),
    .CLK(clknet_leaf_162_wb_clk_i),
    .Q(\soc.ram_step2_read_request ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12171_ (.D(_01199_),
    .CLK(clknet_leaf_161_wb_clk_i),
    .Q(\soc.ram_step1_write_request ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12172_ (.D(_01200_),
    .CLK(clknet_leaf_100_wb_clk_i),
    .Q(\soc.hack_rom_request ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12173_ (.D(_01201_),
    .CLK(clknet_leaf_126_wb_clk_i),
    .Q(\soc.boot_loading_offset[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12174_ (.D(_01202_),
    .CLK(clknet_leaf_126_wb_clk_i),
    .Q(\soc.boot_loading_offset[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12175_ (.D(_01203_),
    .CLK(clknet_leaf_85_wb_clk_i),
    .Q(\soc.boot_loading_offset[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12176_ (.D(_01204_),
    .CLK(clknet_leaf_85_wb_clk_i),
    .Q(\soc.boot_loading_offset[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12177_ (.D(_01205_),
    .CLK(clknet_leaf_85_wb_clk_i),
    .Q(\soc.boot_loading_offset[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _12178_ (.D(_01206_),
    .CLK(clknet_5_15_0_wb_clk_i),
    .Q(\soc.rom_encoder_0.write_enable ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12179_ (.D(_01207_),
    .CLK(clknet_leaf_127_wb_clk_i),
    .Q(\soc.hack_wait_clocks[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12180_ (.D(_01208_),
    .CLK(clknet_leaf_127_wb_clk_i),
    .Q(\soc.hack_wait_clocks[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12181_ (.D(_01209_),
    .CLK(net87),
    .Q(net77));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12182_ (.D(_01210_),
    .CLK(net87),
    .Q(net78));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12183_ (.D(_01211_),
    .CLK(net87),
    .Q(net79));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12184_ (.D(_01212_),
    .CLK(net87),
    .Q(net80));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12185_ (.D(_01213_),
    .CLK(net86),
    .Q(\soc.gpio_i_stored[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12186_ (.D(_01214_),
    .CLK(net87),
    .Q(\soc.gpio_i_stored[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12187_ (.D(_01215_),
    .CLK(net86),
    .Q(\soc.gpio_i_stored[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12188_ (.D(_01216_),
    .CLK(net87),
    .Q(\soc.gpio_i_stored[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12189_ (.D(_01217_),
    .CLK(clknet_leaf_189_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[19][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12190_ (.D(_01218_),
    .CLK(clknet_leaf_219_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[19][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12191_ (.D(_01219_),
    .CLK(clknet_leaf_137_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[19][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12192_ (.D(_01220_),
    .CLK(clknet_leaf_143_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[19][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12193_ (.D(_01221_),
    .CLK(clknet_leaf_139_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[19][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12194_ (.D(_01222_),
    .CLK(clknet_leaf_217_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[19][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12195_ (.D(_01223_),
    .CLK(clknet_leaf_247_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[19][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12196_ (.D(_01224_),
    .CLK(clknet_leaf_194_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[19][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12197_ (.D(_01225_),
    .CLK(clknet_leaf_221_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[19][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12198_ (.D(_01226_),
    .CLK(clknet_leaf_256_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[19][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12199_ (.D(_01227_),
    .CLK(clknet_leaf_20_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[19][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12200_ (.D(_01228_),
    .CLK(clknet_leaf_33_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[19][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12201_ (.D(_01229_),
    .CLK(clknet_leaf_2_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[19][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12202_ (.D(_01230_),
    .CLK(clknet_leaf_40_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[19][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12203_ (.D(_01231_),
    .CLK(clknet_leaf_3_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[19][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12204_ (.D(_01232_),
    .CLK(clknet_leaf_10_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[19][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12205_ (.D(_01233_),
    .CLK(clknet_leaf_79_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[19][16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12206_ (.D(_01234_),
    .CLK(clknet_leaf_79_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[19][17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12207_ (.D(_01235_),
    .CLK(clknet_leaf_76_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[19][18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12208_ (.D(_01236_),
    .CLK(clknet_leaf_67_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[19][19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12209_ (.D(_01237_),
    .CLK(clknet_leaf_51_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[19][20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12210_ (.D(_01238_),
    .CLK(clknet_leaf_241_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[19][21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12211_ (.D(_01239_),
    .CLK(clknet_leaf_252_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[19][22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12212_ (.D(_01240_),
    .CLK(clknet_leaf_234_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[19][23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12213_ (.D(_01241_),
    .CLK(clknet_leaf_305_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[19][24] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12214_ (.D(_01242_),
    .CLK(clknet_leaf_234_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[19][25] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12215_ (.D(_01243_),
    .CLK(clknet_leaf_288_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[19][26] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12216_ (.D(_01244_),
    .CLK(clknet_leaf_264_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[19][27] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12217_ (.D(_01245_),
    .CLK(clknet_leaf_280_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[19][28] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12218_ (.D(_01246_),
    .CLK(clknet_leaf_187_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[29][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12219_ (.D(_01247_),
    .CLK(clknet_leaf_224_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[29][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12220_ (.D(_01248_),
    .CLK(clknet_leaf_262_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[29][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12221_ (.D(_01249_),
    .CLK(clknet_leaf_139_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[29][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12222_ (.D(_01250_),
    .CLK(clknet_leaf_194_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[29][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12223_ (.D(_01251_),
    .CLK(clknet_leaf_176_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[29][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12224_ (.D(_01252_),
    .CLK(clknet_leaf_211_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[29][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12225_ (.D(_01253_),
    .CLK(clknet_leaf_193_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[29][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12226_ (.D(_01254_),
    .CLK(clknet_leaf_177_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[29][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12227_ (.D(_01255_),
    .CLK(clknet_leaf_255_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[29][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12228_ (.D(_01256_),
    .CLK(clknet_leaf_16_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[29][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12229_ (.D(_01257_),
    .CLK(clknet_leaf_36_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[29][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12230_ (.D(_01258_),
    .CLK(clknet_leaf_310_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[29][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12231_ (.D(_01259_),
    .CLK(clknet_leaf_311_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[29][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12232_ (.D(_01260_),
    .CLK(clknet_leaf_316_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[29][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12233_ (.D(_01261_),
    .CLK(clknet_leaf_312_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[29][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12234_ (.D(_01262_),
    .CLK(clknet_leaf_30_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[29][16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12235_ (.D(_01263_),
    .CLK(clknet_leaf_73_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[29][17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12236_ (.D(_01264_),
    .CLK(clknet_leaf_72_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[29][18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12237_ (.D(_01265_),
    .CLK(clknet_leaf_71_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[29][19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12238_ (.D(_01266_),
    .CLK(clknet_leaf_49_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[29][20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12239_ (.D(_01267_),
    .CLK(clknet_leaf_291_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[29][21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12240_ (.D(_01268_),
    .CLK(clknet_leaf_269_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[29][22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12241_ (.D(_01269_),
    .CLK(clknet_leaf_290_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[29][23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12242_ (.D(_01270_),
    .CLK(clknet_leaf_299_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[29][24] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12243_ (.D(_01271_),
    .CLK(clknet_leaf_290_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[29][25] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12244_ (.D(_01272_),
    .CLK(clknet_leaf_294_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[29][26] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12245_ (.D(_01273_),
    .CLK(clknet_leaf_273_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[29][27] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12246_ (.D(_01274_),
    .CLK(clknet_leaf_304_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[29][28] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12247_ (.D(_01275_),
    .CLK(clknet_leaf_187_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[31][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12248_ (.D(_01276_),
    .CLK(clknet_leaf_222_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[31][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12249_ (.D(_01277_),
    .CLK(clknet_leaf_261_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[31][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12250_ (.D(_01278_),
    .CLK(clknet_leaf_135_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[31][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12251_ (.D(_01279_),
    .CLK(clknet_leaf_140_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[31][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12252_ (.D(_01280_),
    .CLK(clknet_leaf_178_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[31][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12253_ (.D(_01281_),
    .CLK(clknet_leaf_210_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[31][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12254_ (.D(_01282_),
    .CLK(clknet_leaf_193_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[31][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12255_ (.D(_01283_),
    .CLK(clknet_leaf_179_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[31][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12256_ (.D(_01284_),
    .CLK(clknet_leaf_257_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[31][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12257_ (.D(_01285_),
    .CLK(clknet_leaf_13_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[31][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12258_ (.D(_01286_),
    .CLK(clknet_leaf_37_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[31][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12259_ (.D(_01287_),
    .CLK(clknet_leaf_311_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[31][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12260_ (.D(_01288_),
    .CLK(clknet_leaf_314_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[31][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12261_ (.D(_01289_),
    .CLK(clknet_leaf_315_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[31][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12262_ (.D(_01290_),
    .CLK(clknet_leaf_311_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[31][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12263_ (.D(_01291_),
    .CLK(clknet_leaf_26_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[31][16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12264_ (.D(_01292_),
    .CLK(clknet_leaf_73_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[31][17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12265_ (.D(_01293_),
    .CLK(clknet_leaf_73_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[31][18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12266_ (.D(_01294_),
    .CLK(clknet_leaf_72_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[31][19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12267_ (.D(_01295_),
    .CLK(clknet_leaf_56_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[31][20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12268_ (.D(_01296_),
    .CLK(clknet_leaf_291_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[31][21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12269_ (.D(_01297_),
    .CLK(clknet_leaf_268_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[31][22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12270_ (.D(_01298_),
    .CLK(clknet_leaf_232_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[31][23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12271_ (.D(_01299_),
    .CLK(clknet_leaf_299_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[31][24] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12272_ (.D(_01300_),
    .CLK(clknet_leaf_231_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[31][25] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12273_ (.D(_01301_),
    .CLK(clknet_leaf_294_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[31][26] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12274_ (.D(_01302_),
    .CLK(clknet_leaf_270_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[31][27] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12275_ (.D(_01303_),
    .CLK(clknet_leaf_303_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[31][28] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12276_ (.D(_01304_),
    .CLK(clknet_leaf_213_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[7][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12277_ (.D(_01305_),
    .CLK(clknet_leaf_245_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[7][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12278_ (.D(_01306_),
    .CLK(clknet_leaf_265_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[7][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12279_ (.D(_01307_),
    .CLK(clknet_leaf_262_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[7][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12280_ (.D(_01308_),
    .CLK(clknet_leaf_258_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[7][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12281_ (.D(_01309_),
    .CLK(clknet_leaf_245_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[7][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12282_ (.D(_01310_),
    .CLK(clknet_leaf_246_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[7][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12283_ (.D(_01311_),
    .CLK(clknet_leaf_244_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[7][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12284_ (.D(_01312_),
    .CLK(clknet_leaf_244_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[7][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12285_ (.D(_01313_),
    .CLK(clknet_leaf_250_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[7][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12286_ (.D(_01314_),
    .CLK(clknet_leaf_13_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[7][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12287_ (.D(_01315_),
    .CLK(clknet_leaf_41_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[7][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12288_ (.D(_01316_),
    .CLK(clknet_leaf_308_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[7][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12289_ (.D(_01317_),
    .CLK(clknet_leaf_312_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[7][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12290_ (.D(_01318_),
    .CLK(clknet_leaf_312_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[7][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12291_ (.D(_01319_),
    .CLK(clknet_leaf_312_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[7][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12292_ (.D(_01320_),
    .CLK(clknet_leaf_75_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[7][16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12293_ (.D(_01321_),
    .CLK(clknet_leaf_80_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[7][17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12294_ (.D(_01322_),
    .CLK(clknet_leaf_80_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[7][18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12295_ (.D(_01323_),
    .CLK(clknet_leaf_73_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[7][19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12296_ (.D(_01324_),
    .CLK(clknet_leaf_49_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[7][20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12297_ (.D(_01325_),
    .CLK(clknet_leaf_292_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[7][21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12298_ (.D(_01326_),
    .CLK(clknet_leaf_268_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[7][22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12299_ (.D(_01327_),
    .CLK(clknet_leaf_286_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[7][23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12300_ (.D(_01328_),
    .CLK(clknet_leaf_300_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[7][24] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12301_ (.D(_01329_),
    .CLK(clknet_leaf_289_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[7][25] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12302_ (.D(_01330_),
    .CLK(clknet_leaf_295_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[7][26] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12303_ (.D(_01331_),
    .CLK(clknet_leaf_272_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[7][27] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12304_ (.D(_01332_),
    .CLK(clknet_leaf_274_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[7][28] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12305_ (.D(_01333_),
    .CLK(clknet_leaf_148_wb_clk_i),
    .Q(\soc.ram_encoder_0.data_out[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12306_ (.D(_01334_),
    .CLK(clknet_leaf_144_wb_clk_i),
    .Q(\soc.ram_encoder_0.data_out[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12307_ (.D(_01335_),
    .CLK(clknet_leaf_144_wb_clk_i),
    .Q(\soc.ram_encoder_0.data_out[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12308_ (.D(_01336_),
    .CLK(clknet_leaf_155_wb_clk_i),
    .Q(\soc.ram_encoder_0.data_out[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12309_ (.D(_01337_),
    .CLK(clknet_leaf_155_wb_clk_i),
    .Q(\soc.ram_encoder_0.data_out[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12310_ (.D(_01338_),
    .CLK(clknet_leaf_154_wb_clk_i),
    .Q(\soc.ram_encoder_0.data_out[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12311_ (.D(_01339_),
    .CLK(clknet_leaf_152_wb_clk_i),
    .Q(\soc.ram_encoder_0.data_out[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12312_ (.D(_01340_),
    .CLK(clknet_leaf_155_wb_clk_i),
    .Q(\soc.ram_encoder_0.data_out[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12313_ (.D(_01341_),
    .CLK(clknet_leaf_155_wb_clk_i),
    .Q(\soc.ram_encoder_0.data_out[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12314_ (.D(_01342_),
    .CLK(clknet_leaf_155_wb_clk_i),
    .Q(\soc.ram_encoder_0.data_out[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12315_ (.D(_01343_),
    .CLK(clknet_leaf_117_wb_clk_i),
    .Q(\soc.ram_encoder_0.data_out[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12316_ (.D(_01344_),
    .CLK(clknet_leaf_117_wb_clk_i),
    .Q(\soc.ram_encoder_0.data_out[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12317_ (.D(_01345_),
    .CLK(clknet_leaf_114_wb_clk_i),
    .Q(\soc.ram_encoder_0.data_out[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12318_ (.D(_01346_),
    .CLK(clknet_leaf_115_wb_clk_i),
    .Q(\soc.ram_encoder_0.data_out[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12319_ (.D(_01347_),
    .CLK(clknet_leaf_115_wb_clk_i),
    .Q(\soc.ram_encoder_0.data_out[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12320_ (.D(_01348_),
    .CLK(clknet_leaf_117_wb_clk_i),
    .Q(\soc.ram_encoder_0.data_out[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12321_ (.D(_01349_),
    .CLK(clknet_leaf_191_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[8][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12322_ (.D(_01350_),
    .CLK(clknet_leaf_222_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[8][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12323_ (.D(_01351_),
    .CLK(clknet_leaf_137_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[8][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12324_ (.D(_01352_),
    .CLK(clknet_leaf_137_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[8][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12325_ (.D(_01353_),
    .CLK(clknet_leaf_197_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[8][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12326_ (.D(_01354_),
    .CLK(clknet_leaf_189_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[8][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12327_ (.D(_01355_),
    .CLK(clknet_leaf_205_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[8][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12328_ (.D(_01356_),
    .CLK(clknet_leaf_193_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[8][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12329_ (.D(_01357_),
    .CLK(clknet_leaf_189_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[8][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12330_ (.D(_01358_),
    .CLK(clknet_leaf_200_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[8][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12331_ (.D(_01359_),
    .CLK(clknet_leaf_13_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[8][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12332_ (.D(_01360_),
    .CLK(clknet_leaf_42_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[8][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12333_ (.D(_01361_),
    .CLK(clknet_leaf_2_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[8][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12334_ (.D(_01362_),
    .CLK(clknet_leaf_7_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[8][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12335_ (.D(_01363_),
    .CLK(clknet_leaf_4_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[8][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12336_ (.D(_01364_),
    .CLK(clknet_leaf_9_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[8][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12337_ (.D(_01365_),
    .CLK(clknet_leaf_26_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[8][16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12338_ (.D(_01366_),
    .CLK(clknet_leaf_24_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[8][17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12339_ (.D(_01367_),
    .CLK(clknet_leaf_26_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[8][18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12340_ (.D(_01368_),
    .CLK(clknet_leaf_31_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[8][19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12341_ (.D(_01369_),
    .CLK(clknet_leaf_53_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[8][20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12342_ (.D(_01370_),
    .CLK(clknet_leaf_283_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[8][21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12343_ (.D(_01371_),
    .CLK(clknet_leaf_252_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[8][22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12344_ (.D(_01372_),
    .CLK(clknet_leaf_238_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[8][23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12345_ (.D(_01373_),
    .CLK(clknet_leaf_306_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[8][24] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12346_ (.D(_01374_),
    .CLK(clknet_leaf_237_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[8][25] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12347_ (.D(_01375_),
    .CLK(clknet_leaf_287_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[8][26] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12348_ (.D(_01376_),
    .CLK(clknet_leaf_271_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[8][27] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12349_ (.D(_01377_),
    .CLK(clknet_leaf_278_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[8][28] ));
 gf180mcu_fd_sc_mcu7t5v0__tieh caravel_hack_soc_225 (.Z(net225));
 gf180mcu_fd_sc_mcu7t5v0__tieh caravel_hack_soc_226 (.Z(net226));
 gf180mcu_fd_sc_mcu7t5v0__tieh caravel_hack_soc_227 (.Z(net227));
 gf180mcu_fd_sc_mcu7t5v0__tieh caravel_hack_soc_228 (.Z(net228));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_0_wb_clk_i (.I(clknet_5_0_0_wb_clk_i),
    .Z(clknet_leaf_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_92 (.ZN(net92));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_93 (.ZN(net93));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_94 (.ZN(net94));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_95 (.ZN(net95));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_96 (.ZN(net96));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_97 (.ZN(net97));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_98 (.ZN(net98));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_99 (.ZN(net99));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_100 (.ZN(net100));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_101 (.ZN(net101));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_102 (.ZN(net102));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_103 (.ZN(net103));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_104 (.ZN(net104));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_105 (.ZN(net105));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_106 (.ZN(net106));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_107 (.ZN(net107));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_108 (.ZN(net108));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_109 (.ZN(net109));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_110 (.ZN(net110));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_111 (.ZN(net111));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_112 (.ZN(net112));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_113 (.ZN(net113));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_114 (.ZN(net114));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_115 (.ZN(net115));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_116 (.ZN(net116));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_117 (.ZN(net117));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_118 (.ZN(net118));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_119 (.ZN(net119));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_120 (.ZN(net120));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_121 (.ZN(net121));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_122 (.ZN(net122));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_123 (.ZN(net123));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_124 (.ZN(net124));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_125 (.ZN(net125));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_126 (.ZN(net126));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_127 (.ZN(net127));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_128 (.ZN(net128));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_129 (.ZN(net129));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_130 (.ZN(net130));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_131 (.ZN(net131));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_132 (.ZN(net132));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_133 (.ZN(net133));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_134 (.ZN(net134));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_135 (.ZN(net135));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_136 (.ZN(net136));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_137 (.ZN(net137));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_138 (.ZN(net138));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_139 (.ZN(net139));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_140 (.ZN(net140));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_141 (.ZN(net141));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_142 (.ZN(net142));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_143 (.ZN(net143));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_144 (.ZN(net144));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_145 (.ZN(net145));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_146 (.ZN(net146));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_147 (.ZN(net147));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_148 (.ZN(net148));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_149 (.ZN(net149));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_150 (.ZN(net150));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_151 (.ZN(net151));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_152 (.ZN(net152));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_153 (.ZN(net153));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_154 (.ZN(net154));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_155 (.ZN(net155));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_156 (.ZN(net156));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_157 (.ZN(net157));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_158 (.ZN(net158));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_159 (.ZN(net159));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_160 (.ZN(net160));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_161 (.ZN(net161));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_162 (.ZN(net162));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_163 (.ZN(net163));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_164 (.ZN(net164));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_165 (.ZN(net165));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_166 (.ZN(net166));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_167 (.ZN(net167));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_168 (.ZN(net168));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_169 (.ZN(net169));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_170 (.ZN(net170));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_171 (.ZN(net171));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_172 (.ZN(net172));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_173 (.ZN(net173));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_174 (.ZN(net174));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_175 (.ZN(net175));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_176 (.ZN(net176));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_177 (.ZN(net177));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_178 (.ZN(net178));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_179 (.ZN(net179));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_180 (.ZN(net180));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_181 (.ZN(net181));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_182 (.ZN(net182));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_183 (.ZN(net183));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_184 (.ZN(net184));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_185 (.ZN(net185));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_186 (.ZN(net186));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_187 (.ZN(net187));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_188 (.ZN(net188));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_189 (.ZN(net189));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_190 (.ZN(net190));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_191 (.ZN(net191));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_192 (.ZN(net192));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_193 (.ZN(net193));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_194 (.ZN(net194));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_195 (.ZN(net195));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_196 (.ZN(net196));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_197 (.ZN(net197));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_198 (.ZN(net198));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_199 (.ZN(net199));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_200 (.ZN(net200));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_201 (.ZN(net201));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_202 (.ZN(net202));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_203 (.ZN(net203));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_204 (.ZN(net204));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_205 (.ZN(net205));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_206 (.ZN(net206));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_207 (.ZN(net207));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_208 (.ZN(net208));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_209 (.ZN(net209));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_210 (.ZN(net210));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_211 (.ZN(net211));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_212 (.ZN(net212));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_213 (.ZN(net213));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_214 (.ZN(net214));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_215 (.ZN(net215));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_216 (.ZN(net216));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_217 (.ZN(net217));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_218 (.ZN(net218));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_219 (.ZN(net219));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_220 (.ZN(net220));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_221 (.ZN(net221));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_222 (.ZN(net222));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_223 (.ZN(net223));
 gf180mcu_fd_sc_mcu7t5v0__tieh caravel_hack_soc_224 (.Z(net224));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12488_ (.I(net49),
    .Z(net46));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12489_ (.I(net49),
    .Z(net47));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12490_ (.I(net49),
    .Z(net48));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12491_ (.I(net53),
    .Z(net50));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12492_ (.I(net53),
    .Z(net51));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12493_ (.I(net53),
    .Z(net52));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12494_ (.I(net57),
    .Z(net54));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12495_ (.I(net57),
    .Z(net55));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12496_ (.I(net57),
    .Z(net56));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_0 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_6 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_7 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_8 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_9 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_10 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_11 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_12 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_13 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_14 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_15 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_16 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_17 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_18 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_19 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_20 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_21 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_22 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_23 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_24 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_25 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_26 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_27 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_28 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_29 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_30 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_31 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_32 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_33 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_34 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_35 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_36 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_37 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_38 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_39 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_40 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_41 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_42 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_43 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_44 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_45 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_46 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_47 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_48 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_49 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_50 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_51 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_52 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_53 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_54 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_55 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_56 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_57 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_58 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_59 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_60 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_61 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_62 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_63 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_64 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_65 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_66 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_67 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_68 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_69 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_70 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_71 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_72 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_73 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_74 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_75 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_76 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_77 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_78 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_79 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_80 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_81 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_82 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_83 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_84 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_85 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_86 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_87 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_88 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_89 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_90 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_91 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_92 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_93 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_94 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_95 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_96 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_97 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_98 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_99 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_100 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_101 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_102 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_103 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_104 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_105 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_106 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_107 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_108 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_109 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_110 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_111 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_112 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_113 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_114 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_115 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_116 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_117 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_118 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_119 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_120 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_121 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_122 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_123 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_124 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_125 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_126 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_127 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_128 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_129 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_130 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_131 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_132 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_133 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_134 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_135 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_136 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_137 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_138 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_139 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_140 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_141 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_142 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_143 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_144 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_145 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_146 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_147 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_148 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_149 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_150 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_151 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_152 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_153 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_154 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_155 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_156 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_157 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_158 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_159 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_160 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_161 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_162 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_163 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_164 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_165 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_166 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_167 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_168 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_169 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_170 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_171 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_172 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_173 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_174 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_175 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_176 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_177 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_178 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_179 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_180 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_181 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_182 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_183 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_184 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_185 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_186 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_187 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_188 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_189 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_190 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_191 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_192 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_193 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_194 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_195 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_196 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_197 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_198 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_199 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_200 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_201 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_202 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_203 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_204 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_205 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_206 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_207 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_208 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_209 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_210 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_211 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_212 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_213 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_214 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_215 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_216 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_217 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_218 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_219 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_220 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_221 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_222 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_223 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_224 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_225 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_226 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_227 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_228 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_229 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_230 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_231 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_232 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_233 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_234 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_235 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_236 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_237 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_238 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_239 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_240 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_241 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_242 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_243 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_244 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_245 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_246 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_247 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_248 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_249 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_250 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_251 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_252 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_253 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_254 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_255 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_256 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_257 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_258 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_259 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_260 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_261 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_262 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_263 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_264 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_265 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_266 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_267 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_268 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_269 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_270 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_271 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_272 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_273 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_274 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_275 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_276 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_277 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_278 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_279 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_280 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_281 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_282 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_283 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_284 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_285 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_286 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_287 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_288 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_289 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_290 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_291 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_292 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_293 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_294 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_295 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_296 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_297 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_298 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_299 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_300 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_301 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_302 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_303 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_304 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_305 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_306 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_307 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_308 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_309 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_310 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_311 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_312 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_313 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_314 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_315 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_316 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_317 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_318 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_319 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_320 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_321 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_322 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_323 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_324 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_325 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_326 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_327 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_328 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_329 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_330 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_331 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_332 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_333 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_334 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_335 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_336 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_337 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_338 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_339 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_340 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_341 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_342 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_343 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_344 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_345 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_346 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_347 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_348 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_349 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_350 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_351 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_352 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_353 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_354 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_355 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_356 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_357 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_358 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_359 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_360 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_361 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_362 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_363 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_364 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_365 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_366 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_367 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_368 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_369 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_370 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_371 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_372 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_373 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_374 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_375 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_376 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_377 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_378 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_379 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_380 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_381 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_382 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_383 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_384 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_385 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_386 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_387 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_388 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_389 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_390 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_391 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_392 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_393 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_394 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_395 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_396 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_397 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_398 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_399 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_400 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_401 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_402 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_403 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_404 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_405 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_406 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_407 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_408 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_409 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_410 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_411 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_412 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_413 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_414 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_415 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_416 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_417 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_418 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_419 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_420 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_421 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_422 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_423 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_424 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_425 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_426 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_427 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_428 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_429 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_430 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_431 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_432 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_433 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_434 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_435 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_436 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_437 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_438 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_439 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_440 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_441 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_442 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_443 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_444 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_445 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_446 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_447 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_448 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_449 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_450 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_451 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_452 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_453 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_454 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_455 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_456 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_457 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_458 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_459 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_460 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_461 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_462 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_463 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_464 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_465 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_466 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_467 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_468 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_469 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_470 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_471 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_472 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_473 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_474 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_475 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_476 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_477 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_478 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_479 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_480 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_481 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_482 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_483 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_484 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_485 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_486 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_487 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_488 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_489 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_490 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_491 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_492 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_4999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_5999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_6595 ();
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1 (.I(io_in[10]),
    .Z(net1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input2 (.I(io_in[11]),
    .Z(net2));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input3 (.I(io_in[12]),
    .Z(net3));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input4 (.I(io_in[13]),
    .Z(net4));
 gf180mcu_fd_sc_mcu7t5v0__dlyd_1 input5 (.I(io_in[16]),
    .Z(net5));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 input6 (.I(io_in[17]),
    .Z(net6));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 input7 (.I(io_in[18]),
    .Z(net7));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input8 (.I(io_in[19]),
    .Z(net8));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input9 (.I(io_in[22]),
    .Z(net9));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input10 (.I(io_in[23]),
    .Z(net10));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input11 (.I(io_in[24]),
    .Z(net11));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input12 (.I(io_in[25]),
    .Z(net12));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 input13 (.I(io_in[26]),
    .Z(net13));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input14 (.I(io_in[30]),
    .Z(net14));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input15 (.I(io_in[31]),
    .Z(net15));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input16 (.I(io_in[32]),
    .Z(net16));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input17 (.I(io_in[33]),
    .Z(net17));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input18 (.I(la_data_in[0]),
    .Z(net18));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input19 (.I(la_data_in[10]),
    .Z(net19));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input20 (.I(la_data_in[11]),
    .Z(net20));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input21 (.I(la_data_in[12]),
    .Z(net21));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input22 (.I(la_data_in[13]),
    .Z(net22));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input23 (.I(la_data_in[14]),
    .Z(net23));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input24 (.I(la_data_in[15]),
    .Z(net24));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input25 (.I(la_data_in[16]),
    .Z(net25));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input26 (.I(la_data_in[17]),
    .Z(net26));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input27 (.I(la_data_in[18]),
    .Z(net27));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input28 (.I(la_data_in[19]),
    .Z(net28));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input29 (.I(la_data_in[1]),
    .Z(net29));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input30 (.I(la_data_in[20]),
    .Z(net30));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input31 (.I(la_data_in[21]),
    .Z(net31));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input32 (.I(la_data_in[22]),
    .Z(net32));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input33 (.I(la_data_in[23]),
    .Z(net33));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input34 (.I(la_data_in[24]),
    .Z(net34));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input35 (.I(la_data_in[25]),
    .Z(net35));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input36 (.I(la_data_in[26]),
    .Z(net36));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input37 (.I(la_data_in[28]),
    .Z(net37));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input38 (.I(la_data_in[2]),
    .Z(net38));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input39 (.I(la_data_in[3]),
    .Z(net39));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input40 (.I(la_data_in[4]),
    .Z(net40));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 input41 (.I(la_data_in[5]),
    .Z(net41));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input42 (.I(la_data_in[6]),
    .Z(net42));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input43 (.I(la_data_in[7]),
    .Z(net43));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input44 (.I(la_data_in[8]),
    .Z(net44));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input45 (.I(la_data_in[9]),
    .Z(net45));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output46 (.I(net46),
    .Z(io_oeb[10]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output47 (.I(net47),
    .Z(io_oeb[11]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output48 (.I(net48),
    .Z(io_oeb[12]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output49 (.I(net49),
    .Z(io_oeb[13]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output50 (.I(net50),
    .Z(io_oeb[16]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output51 (.I(net51),
    .Z(io_oeb[17]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output52 (.I(net52),
    .Z(io_oeb[18]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output53 (.I(net53),
    .Z(io_oeb[19]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output54 (.I(net54),
    .Z(io_oeb[22]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output55 (.I(net55),
    .Z(io_oeb[23]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output56 (.I(net56),
    .Z(io_oeb[24]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output57 (.I(net57),
    .Z(io_oeb[25]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output58 (.I(net58),
    .Z(io_out[10]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output59 (.I(net59),
    .Z(io_out[11]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output60 (.I(net60),
    .Z(io_out[12]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output61 (.I(net61),
    .Z(io_out[13]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output62 (.I(net62),
    .Z(io_out[14]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output63 (.I(net63),
    .Z(io_out[15]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output64 (.I(net64),
    .Z(io_out[16]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output65 (.I(net65),
    .Z(io_out[17]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output66 (.I(net66),
    .Z(io_out[18]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output67 (.I(net67),
    .Z(io_out[19]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output68 (.I(net68),
    .Z(io_out[20]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output69 (.I(net69),
    .Z(io_out[21]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output70 (.I(net70),
    .Z(io_out[22]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output71 (.I(net71),
    .Z(io_out[23]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output72 (.I(net72),
    .Z(io_out[24]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output73 (.I(net73),
    .Z(io_out[25]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output74 (.I(net74),
    .Z(io_out[27]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output75 (.I(net75),
    .Z(io_out[28]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output76 (.I(net76),
    .Z(io_out[29]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output77 (.I(net77),
    .Z(io_out[34]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output78 (.I(net78),
    .Z(io_out[35]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output79 (.I(net79),
    .Z(io_out[36]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output80 (.I(net80),
    .Z(io_out[37]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output81 (.I(net81),
    .Z(io_out[8]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output82 (.I(net82),
    .Z(io_out[9]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output83 (.I(net83),
    .Z(la_data_out[27]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 fanout84 (.I(net85),
    .Z(net84));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 fanout85 (.I(\soc.cpu.AReg.clk ),
    .Z(net85));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 fanout86 (.I(\soc.cpu.AReg.clk ),
    .Z(net86));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 fanout87 (.I(\soc.cpu.AReg.clk ),
    .Z(net87));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 fanout88 (.I(net89),
    .Z(net88));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 fanout89 (.I(net90),
    .Z(net89));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 fanout90 (.I(\soc.cpu.AReg.clk ),
    .Z(net90));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_91 (.ZN(net91));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_1_wb_clk_i (.I(clknet_5_0_0_wb_clk_i),
    .Z(clknet_leaf_1_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_2_wb_clk_i (.I(clknet_5_2_0_wb_clk_i),
    .Z(clknet_leaf_2_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_3_wb_clk_i (.I(clknet_5_2_0_wb_clk_i),
    .Z(clknet_leaf_3_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_4_wb_clk_i (.I(clknet_5_2_0_wb_clk_i),
    .Z(clknet_leaf_4_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_5_wb_clk_i (.I(clknet_5_0_0_wb_clk_i),
    .Z(clknet_leaf_5_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_6_wb_clk_i (.I(clknet_5_0_0_wb_clk_i),
    .Z(clknet_leaf_6_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_7_wb_clk_i (.I(clknet_5_2_0_wb_clk_i),
    .Z(clknet_leaf_7_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_8_wb_clk_i (.I(clknet_5_2_0_wb_clk_i),
    .Z(clknet_leaf_8_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_9_wb_clk_i (.I(clknet_5_3_0_wb_clk_i),
    .Z(clknet_leaf_9_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_10_wb_clk_i (.I(clknet_5_3_0_wb_clk_i),
    .Z(clknet_leaf_10_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_11_wb_clk_i (.I(clknet_5_3_0_wb_clk_i),
    .Z(clknet_leaf_11_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_12_wb_clk_i (.I(clknet_5_2_0_wb_clk_i),
    .Z(clknet_leaf_12_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_13_wb_clk_i (.I(clknet_5_2_0_wb_clk_i),
    .Z(clknet_leaf_13_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_14_wb_clk_i (.I(clknet_5_2_0_wb_clk_i),
    .Z(clknet_leaf_14_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_15_wb_clk_i (.I(clknet_5_2_0_wb_clk_i),
    .Z(clknet_leaf_15_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_16_wb_clk_i (.I(clknet_5_2_0_wb_clk_i),
    .Z(clknet_leaf_16_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_17_wb_clk_i (.I(clknet_5_2_0_wb_clk_i),
    .Z(clknet_leaf_17_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_18_wb_clk_i (.I(clknet_5_2_0_wb_clk_i),
    .Z(clknet_leaf_18_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_19_wb_clk_i (.I(clknet_5_2_0_wb_clk_i),
    .Z(clknet_leaf_19_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_20_wb_clk_i (.I(clknet_5_2_0_wb_clk_i),
    .Z(clknet_leaf_20_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_21_wb_clk_i (.I(clknet_5_8_0_wb_clk_i),
    .Z(clknet_leaf_21_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_22_wb_clk_i (.I(clknet_5_8_0_wb_clk_i),
    .Z(clknet_leaf_22_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_23_wb_clk_i (.I(clknet_5_8_0_wb_clk_i),
    .Z(clknet_leaf_23_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_24_wb_clk_i (.I(clknet_5_8_0_wb_clk_i),
    .Z(clknet_leaf_24_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_25_wb_clk_i (.I(clknet_5_8_0_wb_clk_i),
    .Z(clknet_leaf_25_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_26_wb_clk_i (.I(clknet_5_8_0_wb_clk_i),
    .Z(clknet_leaf_26_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_27_wb_clk_i (.I(clknet_5_8_0_wb_clk_i),
    .Z(clknet_leaf_27_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_28_wb_clk_i (.I(clknet_5_8_0_wb_clk_i),
    .Z(clknet_leaf_28_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_29_wb_clk_i (.I(clknet_5_9_0_wb_clk_i),
    .Z(clknet_leaf_29_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_30_wb_clk_i (.I(clknet_5_9_0_wb_clk_i),
    .Z(clknet_leaf_30_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_31_wb_clk_i (.I(clknet_5_9_0_wb_clk_i),
    .Z(clknet_leaf_31_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_32_wb_clk_i (.I(clknet_5_9_0_wb_clk_i),
    .Z(clknet_leaf_32_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_33_wb_clk_i (.I(clknet_5_9_0_wb_clk_i),
    .Z(clknet_leaf_33_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_34_wb_clk_i (.I(clknet_5_9_0_wb_clk_i),
    .Z(clknet_leaf_34_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_35_wb_clk_i (.I(clknet_5_9_0_wb_clk_i),
    .Z(clknet_leaf_35_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_36_wb_clk_i (.I(clknet_5_2_0_wb_clk_i),
    .Z(clknet_leaf_36_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_37_wb_clk_i (.I(clknet_5_3_0_wb_clk_i),
    .Z(clknet_leaf_37_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_38_wb_clk_i (.I(clknet_5_3_0_wb_clk_i),
    .Z(clknet_leaf_38_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_39_wb_clk_i (.I(clknet_5_3_0_wb_clk_i),
    .Z(clknet_leaf_39_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_40_wb_clk_i (.I(clknet_5_3_0_wb_clk_i),
    .Z(clknet_leaf_40_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_41_wb_clk_i (.I(clknet_5_6_0_wb_clk_i),
    .Z(clknet_leaf_41_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_42_wb_clk_i (.I(clknet_5_3_0_wb_clk_i),
    .Z(clknet_leaf_42_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_43_wb_clk_i (.I(clknet_5_6_0_wb_clk_i),
    .Z(clknet_leaf_43_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_44_wb_clk_i (.I(clknet_5_6_0_wb_clk_i),
    .Z(clknet_leaf_44_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_45_wb_clk_i (.I(clknet_5_6_0_wb_clk_i),
    .Z(clknet_leaf_45_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_46_wb_clk_i (.I(clknet_5_3_0_wb_clk_i),
    .Z(clknet_leaf_46_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_47_wb_clk_i (.I(clknet_5_9_0_wb_clk_i),
    .Z(clknet_leaf_47_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_48_wb_clk_i (.I(clknet_5_12_0_wb_clk_i),
    .Z(clknet_leaf_48_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_49_wb_clk_i (.I(clknet_5_13_0_wb_clk_i),
    .Z(clknet_leaf_49_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_50_wb_clk_i (.I(clknet_5_6_0_wb_clk_i),
    .Z(clknet_leaf_50_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_51_wb_clk_i (.I(clknet_5_6_0_wb_clk_i),
    .Z(clknet_leaf_51_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_52_wb_clk_i (.I(clknet_5_13_0_wb_clk_i),
    .Z(clknet_leaf_52_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_53_wb_clk_i (.I(clknet_5_13_0_wb_clk_i),
    .Z(clknet_leaf_53_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_54_wb_clk_i (.I(clknet_5_24_0_wb_clk_i),
    .Z(clknet_leaf_54_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_55_wb_clk_i (.I(clknet_5_24_0_wb_clk_i),
    .Z(clknet_leaf_55_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_56_wb_clk_i (.I(clknet_5_13_0_wb_clk_i),
    .Z(clknet_leaf_56_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_58_wb_clk_i (.I(clknet_5_12_0_wb_clk_i),
    .Z(clknet_leaf_58_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_59_wb_clk_i (.I(clknet_5_13_0_wb_clk_i),
    .Z(clknet_leaf_59_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_60_wb_clk_i (.I(clknet_5_12_0_wb_clk_i),
    .Z(clknet_leaf_60_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_61_wb_clk_i (.I(clknet_5_9_0_wb_clk_i),
    .Z(clknet_leaf_61_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_62_wb_clk_i (.I(clknet_5_12_0_wb_clk_i),
    .Z(clknet_leaf_62_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_63_wb_clk_i (.I(clknet_5_12_0_wb_clk_i),
    .Z(clknet_leaf_63_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_64_wb_clk_i (.I(clknet_5_12_0_wb_clk_i),
    .Z(clknet_leaf_64_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_65_wb_clk_i (.I(clknet_5_11_0_wb_clk_i),
    .Z(clknet_leaf_65_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_66_wb_clk_i (.I(clknet_5_11_0_wb_clk_i),
    .Z(clknet_leaf_66_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_67_wb_clk_i (.I(clknet_5_11_0_wb_clk_i),
    .Z(clknet_leaf_67_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_68_wb_clk_i (.I(clknet_5_11_0_wb_clk_i),
    .Z(clknet_leaf_68_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_69_wb_clk_i (.I(clknet_5_11_0_wb_clk_i),
    .Z(clknet_leaf_69_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_70_wb_clk_i (.I(clknet_5_9_0_wb_clk_i),
    .Z(clknet_leaf_70_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_71_wb_clk_i (.I(clknet_5_9_0_wb_clk_i),
    .Z(clknet_leaf_71_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_72_wb_clk_i (.I(clknet_5_9_0_wb_clk_i),
    .Z(clknet_leaf_72_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_73_wb_clk_i (.I(clknet_5_8_0_wb_clk_i),
    .Z(clknet_leaf_73_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_74_wb_clk_i (.I(clknet_5_9_0_wb_clk_i),
    .Z(clknet_leaf_74_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_75_wb_clk_i (.I(clknet_5_8_0_wb_clk_i),
    .Z(clknet_leaf_75_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_76_wb_clk_i (.I(clknet_5_8_0_wb_clk_i),
    .Z(clknet_leaf_76_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_77_wb_clk_i (.I(clknet_5_8_0_wb_clk_i),
    .Z(clknet_leaf_77_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_78_wb_clk_i (.I(clknet_5_8_0_wb_clk_i),
    .Z(clknet_leaf_78_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_79_wb_clk_i (.I(clknet_5_10_0_wb_clk_i),
    .Z(clknet_leaf_79_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_80_wb_clk_i (.I(clknet_5_10_0_wb_clk_i),
    .Z(clknet_leaf_80_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_81_wb_clk_i (.I(clknet_5_10_0_wb_clk_i),
    .Z(clknet_leaf_81_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_82_wb_clk_i (.I(clknet_5_10_0_wb_clk_i),
    .Z(clknet_leaf_82_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_83_wb_clk_i (.I(clknet_5_10_0_wb_clk_i),
    .Z(clknet_leaf_83_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_85_wb_clk_i (.I(clknet_5_14_0_wb_clk_i),
    .Z(clknet_leaf_85_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_86_wb_clk_i (.I(clknet_5_14_0_wb_clk_i),
    .Z(clknet_leaf_86_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_87_wb_clk_i (.I(clknet_5_11_0_wb_clk_i),
    .Z(clknet_leaf_87_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_89_wb_clk_i (.I(clknet_5_10_0_wb_clk_i),
    .Z(clknet_leaf_89_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_92_wb_clk_i (.I(clknet_5_14_0_wb_clk_i),
    .Z(clknet_leaf_92_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_93_wb_clk_i (.I(clknet_5_14_0_wb_clk_i),
    .Z(clknet_leaf_93_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_95_wb_clk_i (.I(clknet_5_11_0_wb_clk_i),
    .Z(clknet_leaf_95_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_96_wb_clk_i (.I(clknet_5_11_0_wb_clk_i),
    .Z(clknet_leaf_96_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_97_wb_clk_i (.I(clknet_5_14_0_wb_clk_i),
    .Z(clknet_leaf_97_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_98_wb_clk_i (.I(clknet_5_14_0_wb_clk_i),
    .Z(clknet_leaf_98_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_99_wb_clk_i (.I(clknet_5_14_0_wb_clk_i),
    .Z(clknet_leaf_99_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_100_wb_clk_i (.I(clknet_5_14_0_wb_clk_i),
    .Z(clknet_leaf_100_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_101_wb_clk_i (.I(clknet_5_14_0_wb_clk_i),
    .Z(clknet_leaf_101_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_102_wb_clk_i (.I(clknet_5_15_0_wb_clk_i),
    .Z(clknet_leaf_102_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_104_wb_clk_i (.I(clknet_5_14_0_wb_clk_i),
    .Z(clknet_leaf_104_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_105_wb_clk_i (.I(clknet_5_14_0_wb_clk_i),
    .Z(clknet_leaf_105_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_106_wb_clk_i (.I(clknet_5_14_0_wb_clk_i),
    .Z(clknet_leaf_106_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_107_wb_clk_i (.I(clknet_5_15_0_wb_clk_i),
    .Z(clknet_leaf_107_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_108_wb_clk_i (.I(clknet_5_15_0_wb_clk_i),
    .Z(clknet_leaf_108_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_109_wb_clk_i (.I(clknet_5_15_0_wb_clk_i),
    .Z(clknet_leaf_109_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_110_wb_clk_i (.I(clknet_5_15_0_wb_clk_i),
    .Z(clknet_leaf_110_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_111_wb_clk_i (.I(clknet_opt_3_0_wb_clk_i),
    .Z(clknet_leaf_111_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_112_wb_clk_i (.I(clknet_opt_4_0_wb_clk_i),
    .Z(clknet_leaf_112_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_113_wb_clk_i (.I(clknet_5_26_0_wb_clk_i),
    .Z(clknet_leaf_113_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_114_wb_clk_i (.I(clknet_5_26_0_wb_clk_i),
    .Z(clknet_leaf_114_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_115_wb_clk_i (.I(clknet_5_26_0_wb_clk_i),
    .Z(clknet_leaf_115_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_117_wb_clk_i (.I(clknet_5_26_0_wb_clk_i),
    .Z(clknet_leaf_117_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_118_wb_clk_i (.I(clknet_5_26_0_wb_clk_i),
    .Z(clknet_leaf_118_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_119_wb_clk_i (.I(clknet_5_26_0_wb_clk_i),
    .Z(clknet_leaf_119_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_121_wb_clk_i (.I(clknet_5_15_0_wb_clk_i),
    .Z(clknet_leaf_121_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_122_wb_clk_i (.I(clknet_5_15_0_wb_clk_i),
    .Z(clknet_leaf_122_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_123_wb_clk_i (.I(clknet_5_15_0_wb_clk_i),
    .Z(clknet_leaf_123_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_124_wb_clk_i (.I(clknet_5_13_0_wb_clk_i),
    .Z(clknet_leaf_124_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_125_wb_clk_i (.I(clknet_5_12_0_wb_clk_i),
    .Z(clknet_leaf_125_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_126_wb_clk_i (.I(clknet_5_14_0_wb_clk_i),
    .Z(clknet_leaf_126_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_127_wb_clk_i (.I(clknet_5_13_0_wb_clk_i),
    .Z(clknet_leaf_127_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_128_wb_clk_i (.I(clknet_5_13_0_wb_clk_i),
    .Z(clknet_leaf_128_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_129_wb_clk_i (.I(clknet_5_12_0_wb_clk_i),
    .Z(clknet_leaf_129_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_130_wb_clk_i (.I(clknet_5_13_0_wb_clk_i),
    .Z(clknet_leaf_130_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_132_wb_clk_i (.I(clknet_5_24_0_wb_clk_i),
    .Z(clknet_leaf_132_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_134_wb_clk_i (.I(clknet_5_24_0_wb_clk_i),
    .Z(clknet_leaf_134_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_135_wb_clk_i (.I(clknet_5_24_0_wb_clk_i),
    .Z(clknet_leaf_135_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_136_wb_clk_i (.I(clknet_5_24_0_wb_clk_i),
    .Z(clknet_leaf_136_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_137_wb_clk_i (.I(clknet_5_24_0_wb_clk_i),
    .Z(clknet_leaf_137_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_138_wb_clk_i (.I(clknet_5_25_0_wb_clk_i),
    .Z(clknet_leaf_138_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_139_wb_clk_i (.I(clknet_5_24_0_wb_clk_i),
    .Z(clknet_leaf_139_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_140_wb_clk_i (.I(clknet_5_25_0_wb_clk_i),
    .Z(clknet_leaf_140_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_141_wb_clk_i (.I(clknet_5_25_0_wb_clk_i),
    .Z(clknet_leaf_141_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_142_wb_clk_i (.I(clknet_5_25_0_wb_clk_i),
    .Z(clknet_leaf_142_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_143_wb_clk_i (.I(clknet_5_24_0_wb_clk_i),
    .Z(clknet_leaf_143_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_144_wb_clk_i (.I(clknet_5_28_0_wb_clk_i),
    .Z(clknet_leaf_144_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_145_wb_clk_i (.I(clknet_5_25_0_wb_clk_i),
    .Z(clknet_leaf_145_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_146_wb_clk_i (.I(clknet_5_28_0_wb_clk_i),
    .Z(clknet_leaf_146_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_147_wb_clk_i (.I(clknet_5_28_0_wb_clk_i),
    .Z(clknet_leaf_147_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_148_wb_clk_i (.I(clknet_5_28_0_wb_clk_i),
    .Z(clknet_leaf_148_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_149_wb_clk_i (.I(clknet_5_29_0_wb_clk_i),
    .Z(clknet_leaf_149_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_150_wb_clk_i (.I(clknet_5_31_0_wb_clk_i),
    .Z(clknet_leaf_150_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_151_wb_clk_i (.I(clknet_5_30_0_wb_clk_i),
    .Z(clknet_leaf_151_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_152_wb_clk_i (.I(clknet_5_30_0_wb_clk_i),
    .Z(clknet_leaf_152_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_153_wb_clk_i (.I(clknet_5_30_0_wb_clk_i),
    .Z(clknet_leaf_153_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_154_wb_clk_i (.I(clknet_5_30_0_wb_clk_i),
    .Z(clknet_leaf_154_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_155_wb_clk_i (.I(clknet_5_30_0_wb_clk_i),
    .Z(clknet_leaf_155_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_156_wb_clk_i (.I(clknet_5_30_0_wb_clk_i),
    .Z(clknet_leaf_156_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_157_wb_clk_i (.I(clknet_5_27_0_wb_clk_i),
    .Z(clknet_leaf_157_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_158_wb_clk_i (.I(clknet_5_27_0_wb_clk_i),
    .Z(clknet_leaf_158_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_159_wb_clk_i (.I(clknet_5_27_0_wb_clk_i),
    .Z(clknet_leaf_159_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_160_wb_clk_i (.I(clknet_5_27_0_wb_clk_i),
    .Z(clknet_leaf_160_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_161_wb_clk_i (.I(clknet_5_27_0_wb_clk_i),
    .Z(clknet_leaf_161_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_162_wb_clk_i (.I(clknet_5_27_0_wb_clk_i),
    .Z(clknet_leaf_162_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_163_wb_clk_i (.I(clknet_5_27_0_wb_clk_i),
    .Z(clknet_leaf_163_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_164_wb_clk_i (.I(clknet_5_27_0_wb_clk_i),
    .Z(clknet_leaf_164_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_165_wb_clk_i (.I(clknet_5_30_0_wb_clk_i),
    .Z(clknet_leaf_165_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_166_wb_clk_i (.I(clknet_5_30_0_wb_clk_i),
    .Z(clknet_leaf_166_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_167_wb_clk_i (.I(clknet_5_30_0_wb_clk_i),
    .Z(clknet_leaf_167_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_168_wb_clk_i (.I(clknet_5_30_0_wb_clk_i),
    .Z(clknet_leaf_168_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_169_wb_clk_i (.I(clknet_5_31_0_wb_clk_i),
    .Z(clknet_leaf_169_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_170_wb_clk_i (.I(clknet_5_31_0_wb_clk_i),
    .Z(clknet_leaf_170_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_173_wb_clk_i (.I(clknet_opt_5_0_wb_clk_i),
    .Z(clknet_leaf_173_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_175_wb_clk_i (.I(clknet_5_23_0_wb_clk_i),
    .Z(clknet_leaf_175_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_176_wb_clk_i (.I(clknet_5_23_0_wb_clk_i),
    .Z(clknet_leaf_176_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_177_wb_clk_i (.I(clknet_5_23_0_wb_clk_i),
    .Z(clknet_leaf_177_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_178_wb_clk_i (.I(clknet_5_23_0_wb_clk_i),
    .Z(clknet_leaf_178_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_179_wb_clk_i (.I(clknet_5_23_0_wb_clk_i),
    .Z(clknet_leaf_179_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_180_wb_clk_i (.I(clknet_5_29_0_wb_clk_i),
    .Z(clknet_leaf_180_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_183_wb_clk_i (.I(clknet_5_29_0_wb_clk_i),
    .Z(clknet_leaf_183_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_184_wb_clk_i (.I(clknet_5_29_0_wb_clk_i),
    .Z(clknet_leaf_184_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_185_wb_clk_i (.I(clknet_5_28_0_wb_clk_i),
    .Z(clknet_leaf_185_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_186_wb_clk_i (.I(clknet_5_28_0_wb_clk_i),
    .Z(clknet_leaf_186_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_187_wb_clk_i (.I(clknet_5_29_0_wb_clk_i),
    .Z(clknet_leaf_187_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_188_wb_clk_i (.I(clknet_5_29_0_wb_clk_i),
    .Z(clknet_leaf_188_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_189_wb_clk_i (.I(clknet_5_22_0_wb_clk_i),
    .Z(clknet_leaf_189_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_190_wb_clk_i (.I(clknet_5_22_0_wb_clk_i),
    .Z(clknet_leaf_190_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_191_wb_clk_i (.I(clknet_5_22_0_wb_clk_i),
    .Z(clknet_leaf_191_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_192_wb_clk_i (.I(clknet_5_28_0_wb_clk_i),
    .Z(clknet_leaf_192_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_193_wb_clk_i (.I(clknet_5_28_0_wb_clk_i),
    .Z(clknet_leaf_193_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_194_wb_clk_i (.I(clknet_5_25_0_wb_clk_i),
    .Z(clknet_leaf_194_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_195_wb_clk_i (.I(clknet_5_25_0_wb_clk_i),
    .Z(clknet_leaf_195_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_196_wb_clk_i (.I(clknet_5_25_0_wb_clk_i),
    .Z(clknet_leaf_196_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_197_wb_clk_i (.I(clknet_5_25_0_wb_clk_i),
    .Z(clknet_leaf_197_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_198_wb_clk_i (.I(clknet_5_25_0_wb_clk_i),
    .Z(clknet_leaf_198_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_199_wb_clk_i (.I(clknet_5_18_0_wb_clk_i),
    .Z(clknet_leaf_199_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_200_wb_clk_i (.I(clknet_5_19_0_wb_clk_i),
    .Z(clknet_leaf_200_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_201_wb_clk_i (.I(clknet_5_19_0_wb_clk_i),
    .Z(clknet_leaf_201_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_202_wb_clk_i (.I(clknet_5_19_0_wb_clk_i),
    .Z(clknet_leaf_202_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_203_wb_clk_i (.I(clknet_5_22_0_wb_clk_i),
    .Z(clknet_leaf_203_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_205_wb_clk_i (.I(clknet_5_22_0_wb_clk_i),
    .Z(clknet_leaf_205_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_207_wb_clk_i (.I(clknet_5_22_0_wb_clk_i),
    .Z(clknet_leaf_207_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_208_wb_clk_i (.I(clknet_5_22_0_wb_clk_i),
    .Z(clknet_leaf_208_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_210_wb_clk_i (.I(clknet_5_20_0_wb_clk_i),
    .Z(clknet_leaf_210_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_211_wb_clk_i (.I(clknet_5_20_0_wb_clk_i),
    .Z(clknet_leaf_211_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_212_wb_clk_i (.I(clknet_5_20_0_wb_clk_i),
    .Z(clknet_leaf_212_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_213_wb_clk_i (.I(clknet_5_20_0_wb_clk_i),
    .Z(clknet_leaf_213_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_214_wb_clk_i (.I(clknet_5_20_0_wb_clk_i),
    .Z(clknet_leaf_214_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_215_wb_clk_i (.I(clknet_5_21_0_wb_clk_i),
    .Z(clknet_leaf_215_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_216_wb_clk_i (.I(clknet_5_21_0_wb_clk_i),
    .Z(clknet_leaf_216_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_217_wb_clk_i (.I(clknet_5_21_0_wb_clk_i),
    .Z(clknet_leaf_217_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_218_wb_clk_i (.I(clknet_5_21_0_wb_clk_i),
    .Z(clknet_leaf_218_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_219_wb_clk_i (.I(clknet_5_21_0_wb_clk_i),
    .Z(clknet_leaf_219_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_220_wb_clk_i (.I(clknet_5_21_0_wb_clk_i),
    .Z(clknet_leaf_220_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_221_wb_clk_i (.I(clknet_5_23_0_wb_clk_i),
    .Z(clknet_leaf_221_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_222_wb_clk_i (.I(clknet_5_23_0_wb_clk_i),
    .Z(clknet_leaf_222_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_224_wb_clk_i (.I(clknet_5_23_0_wb_clk_i),
    .Z(clknet_leaf_224_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_226_wb_clk_i (.I(clknet_5_21_0_wb_clk_i),
    .Z(clknet_leaf_226_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_227_wb_clk_i (.I(clknet_5_20_0_wb_clk_i),
    .Z(clknet_leaf_227_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_228_wb_clk_i (.I(clknet_5_20_0_wb_clk_i),
    .Z(clknet_leaf_228_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_229_wb_clk_i (.I(clknet_5_16_0_wb_clk_i),
    .Z(clknet_leaf_229_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_230_wb_clk_i (.I(clknet_5_16_0_wb_clk_i),
    .Z(clknet_leaf_230_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_231_wb_clk_i (.I(clknet_5_5_0_wb_clk_i),
    .Z(clknet_leaf_231_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_232_wb_clk_i (.I(clknet_5_5_0_wb_clk_i),
    .Z(clknet_leaf_232_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_233_wb_clk_i (.I(clknet_5_5_0_wb_clk_i),
    .Z(clknet_leaf_233_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_234_wb_clk_i (.I(clknet_5_16_0_wb_clk_i),
    .Z(clknet_leaf_234_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_235_wb_clk_i (.I(clknet_5_16_0_wb_clk_i),
    .Z(clknet_leaf_235_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_236_wb_clk_i (.I(clknet_5_5_0_wb_clk_i),
    .Z(clknet_leaf_236_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_237_wb_clk_i (.I(clknet_5_5_0_wb_clk_i),
    .Z(clknet_leaf_237_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_238_wb_clk_i (.I(clknet_5_7_0_wb_clk_i),
    .Z(clknet_leaf_238_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_239_wb_clk_i (.I(clknet_5_16_0_wb_clk_i),
    .Z(clknet_leaf_239_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_240_wb_clk_i (.I(clknet_5_17_0_wb_clk_i),
    .Z(clknet_leaf_240_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_241_wb_clk_i (.I(clknet_5_16_0_wb_clk_i),
    .Z(clknet_leaf_241_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_242_wb_clk_i (.I(clknet_5_16_0_wb_clk_i),
    .Z(clknet_leaf_242_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_243_wb_clk_i (.I(clknet_5_17_0_wb_clk_i),
    .Z(clknet_leaf_243_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_244_wb_clk_i (.I(clknet_5_17_0_wb_clk_i),
    .Z(clknet_leaf_244_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_245_wb_clk_i (.I(clknet_5_17_0_wb_clk_i),
    .Z(clknet_leaf_245_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_246_wb_clk_i (.I(clknet_5_17_0_wb_clk_i),
    .Z(clknet_leaf_246_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_247_wb_clk_i (.I(clknet_5_19_0_wb_clk_i),
    .Z(clknet_leaf_247_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_248_wb_clk_i (.I(clknet_5_19_0_wb_clk_i),
    .Z(clknet_leaf_248_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_249_wb_clk_i (.I(clknet_5_17_0_wb_clk_i),
    .Z(clknet_leaf_249_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_250_wb_clk_i (.I(clknet_5_17_0_wb_clk_i),
    .Z(clknet_leaf_250_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_251_wb_clk_i (.I(clknet_5_7_0_wb_clk_i),
    .Z(clknet_leaf_251_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_252_wb_clk_i (.I(clknet_5_7_0_wb_clk_i),
    .Z(clknet_leaf_252_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_253_wb_clk_i (.I(clknet_5_7_0_wb_clk_i),
    .Z(clknet_leaf_253_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_254_wb_clk_i (.I(clknet_5_7_0_wb_clk_i),
    .Z(clknet_leaf_254_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_255_wb_clk_i (.I(clknet_5_18_0_wb_clk_i),
    .Z(clknet_leaf_255_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_256_wb_clk_i (.I(clknet_5_18_0_wb_clk_i),
    .Z(clknet_leaf_256_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_257_wb_clk_i (.I(clknet_5_18_0_wb_clk_i),
    .Z(clknet_leaf_257_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_258_wb_clk_i (.I(clknet_5_18_0_wb_clk_i),
    .Z(clknet_leaf_258_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_259_wb_clk_i (.I(clknet_5_18_0_wb_clk_i),
    .Z(clknet_leaf_259_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_260_wb_clk_i (.I(clknet_5_18_0_wb_clk_i),
    .Z(clknet_leaf_260_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_261_wb_clk_i (.I(clknet_5_7_0_wb_clk_i),
    .Z(clknet_leaf_261_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_262_wb_clk_i (.I(clknet_5_7_0_wb_clk_i),
    .Z(clknet_leaf_262_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_263_wb_clk_i (.I(clknet_5_7_0_wb_clk_i),
    .Z(clknet_leaf_263_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_264_wb_clk_i (.I(clknet_5_6_0_wb_clk_i),
    .Z(clknet_leaf_264_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_265_wb_clk_i (.I(clknet_5_7_0_wb_clk_i),
    .Z(clknet_leaf_265_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_266_wb_clk_i (.I(clknet_5_7_0_wb_clk_i),
    .Z(clknet_leaf_266_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_267_wb_clk_i (.I(clknet_5_7_0_wb_clk_i),
    .Z(clknet_leaf_267_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_268_wb_clk_i (.I(clknet_5_7_0_wb_clk_i),
    .Z(clknet_leaf_268_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_269_wb_clk_i (.I(clknet_5_7_0_wb_clk_i),
    .Z(clknet_leaf_269_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_270_wb_clk_i (.I(clknet_5_6_0_wb_clk_i),
    .Z(clknet_leaf_270_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_271_wb_clk_i (.I(clknet_5_6_0_wb_clk_i),
    .Z(clknet_leaf_271_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_272_wb_clk_i (.I(clknet_5_6_0_wb_clk_i),
    .Z(clknet_leaf_272_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_273_wb_clk_i (.I(clknet_5_6_0_wb_clk_i),
    .Z(clknet_leaf_273_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_274_wb_clk_i (.I(clknet_5_6_0_wb_clk_i),
    .Z(clknet_leaf_274_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_276_wb_clk_i (.I(clknet_5_6_0_wb_clk_i),
    .Z(clknet_leaf_276_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_277_wb_clk_i (.I(clknet_5_4_0_wb_clk_i),
    .Z(clknet_leaf_277_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_278_wb_clk_i (.I(clknet_5_4_0_wb_clk_i),
    .Z(clknet_leaf_278_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_279_wb_clk_i (.I(clknet_5_4_0_wb_clk_i),
    .Z(clknet_leaf_279_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_280_wb_clk_i (.I(clknet_5_4_0_wb_clk_i),
    .Z(clknet_leaf_280_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_281_wb_clk_i (.I(clknet_5_4_0_wb_clk_i),
    .Z(clknet_leaf_281_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_282_wb_clk_i (.I(clknet_5_7_0_wb_clk_i),
    .Z(clknet_leaf_282_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_283_wb_clk_i (.I(clknet_5_7_0_wb_clk_i),
    .Z(clknet_leaf_283_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_284_wb_clk_i (.I(clknet_5_7_0_wb_clk_i),
    .Z(clknet_leaf_284_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_285_wb_clk_i (.I(clknet_5_5_0_wb_clk_i),
    .Z(clknet_leaf_285_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_286_wb_clk_i (.I(clknet_5_5_0_wb_clk_i),
    .Z(clknet_leaf_286_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_287_wb_clk_i (.I(clknet_5_5_0_wb_clk_i),
    .Z(clknet_leaf_287_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_288_wb_clk_i (.I(clknet_5_4_0_wb_clk_i),
    .Z(clknet_leaf_288_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_289_wb_clk_i (.I(clknet_5_5_0_wb_clk_i),
    .Z(clknet_leaf_289_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_290_wb_clk_i (.I(clknet_5_5_0_wb_clk_i),
    .Z(clknet_leaf_290_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_291_wb_clk_i (.I(clknet_5_5_0_wb_clk_i),
    .Z(clknet_leaf_291_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_292_wb_clk_i (.I(clknet_5_5_0_wb_clk_i),
    .Z(clknet_leaf_292_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_293_wb_clk_i (.I(clknet_5_4_0_wb_clk_i),
    .Z(clknet_leaf_293_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_294_wb_clk_i (.I(clknet_5_4_0_wb_clk_i),
    .Z(clknet_leaf_294_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_295_wb_clk_i (.I(clknet_5_4_0_wb_clk_i),
    .Z(clknet_leaf_295_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_296_wb_clk_i (.I(clknet_5_4_0_wb_clk_i),
    .Z(clknet_leaf_296_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_297_wb_clk_i (.I(clknet_5_4_0_wb_clk_i),
    .Z(clknet_leaf_297_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_298_wb_clk_i (.I(clknet_5_1_0_wb_clk_i),
    .Z(clknet_leaf_298_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_299_wb_clk_i (.I(clknet_5_1_0_wb_clk_i),
    .Z(clknet_leaf_299_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_300_wb_clk_i (.I(clknet_5_1_0_wb_clk_i),
    .Z(clknet_leaf_300_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_301_wb_clk_i (.I(clknet_5_1_0_wb_clk_i),
    .Z(clknet_leaf_301_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_302_wb_clk_i (.I(clknet_5_4_0_wb_clk_i),
    .Z(clknet_leaf_302_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_303_wb_clk_i (.I(clknet_5_4_0_wb_clk_i),
    .Z(clknet_leaf_303_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_304_wb_clk_i (.I(clknet_5_1_0_wb_clk_i),
    .Z(clknet_leaf_304_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_305_wb_clk_i (.I(clknet_5_1_0_wb_clk_i),
    .Z(clknet_leaf_305_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_306_wb_clk_i (.I(clknet_5_3_0_wb_clk_i),
    .Z(clknet_leaf_306_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_307_wb_clk_i (.I(clknet_5_3_0_wb_clk_i),
    .Z(clknet_leaf_307_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_308_wb_clk_i (.I(clknet_5_1_0_wb_clk_i),
    .Z(clknet_leaf_308_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_309_wb_clk_i (.I(clknet_5_1_0_wb_clk_i),
    .Z(clknet_leaf_309_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_310_wb_clk_i (.I(clknet_5_0_0_wb_clk_i),
    .Z(clknet_leaf_310_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_311_wb_clk_i (.I(clknet_5_1_0_wb_clk_i),
    .Z(clknet_leaf_311_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_312_wb_clk_i (.I(clknet_5_1_0_wb_clk_i),
    .Z(clknet_leaf_312_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_313_wb_clk_i (.I(clknet_5_1_0_wb_clk_i),
    .Z(clknet_leaf_313_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_314_wb_clk_i (.I(clknet_5_1_0_wb_clk_i),
    .Z(clknet_leaf_314_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_315_wb_clk_i (.I(clknet_5_0_0_wb_clk_i),
    .Z(clknet_leaf_315_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_316_wb_clk_i (.I(clknet_5_0_0_wb_clk_i),
    .Z(clknet_leaf_316_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_317_wb_clk_i (.I(clknet_5_0_0_wb_clk_i),
    .Z(clknet_leaf_317_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_318_wb_clk_i (.I(clknet_5_0_0_wb_clk_i),
    .Z(clknet_leaf_318_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_319_wb_clk_i (.I(clknet_5_0_0_wb_clk_i),
    .Z(clknet_leaf_319_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_320_wb_clk_i (.I(clknet_5_0_0_wb_clk_i),
    .Z(clknet_leaf_320_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_321_wb_clk_i (.I(clknet_5_0_0_wb_clk_i),
    .Z(clknet_leaf_321_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_0_wb_clk_i (.I(wb_clk_i),
    .Z(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_2_0_0_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_2_0_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_2_1_0_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_2_1_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_2_2_0_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_2_2_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_2_3_0_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_2_3_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_0_0_wb_clk_i (.I(clknet_2_0_0_wb_clk_i),
    .Z(clknet_3_0_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_1_0_wb_clk_i (.I(clknet_2_0_0_wb_clk_i),
    .Z(clknet_3_1_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_2_0_wb_clk_i (.I(clknet_2_1_0_wb_clk_i),
    .Z(clknet_3_2_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_3_0_wb_clk_i (.I(clknet_2_1_0_wb_clk_i),
    .Z(clknet_3_3_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_4_0_wb_clk_i (.I(clknet_2_2_0_wb_clk_i),
    .Z(clknet_3_4_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_5_0_wb_clk_i (.I(clknet_2_2_0_wb_clk_i),
    .Z(clknet_3_5_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_6_0_wb_clk_i (.I(clknet_2_3_0_wb_clk_i),
    .Z(clknet_3_6_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_7_0_wb_clk_i (.I(clknet_2_3_0_wb_clk_i),
    .Z(clknet_3_7_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_4_0_0_wb_clk_i (.I(clknet_3_0_0_wb_clk_i),
    .Z(clknet_4_0_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_4_1_0_wb_clk_i (.I(clknet_3_0_0_wb_clk_i),
    .Z(clknet_4_1_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_4_2_0_wb_clk_i (.I(clknet_3_1_0_wb_clk_i),
    .Z(clknet_4_2_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_4_3_0_wb_clk_i (.I(clknet_3_1_0_wb_clk_i),
    .Z(clknet_4_3_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_4_4_0_wb_clk_i (.I(clknet_3_2_0_wb_clk_i),
    .Z(clknet_4_4_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_4_5_0_wb_clk_i (.I(clknet_3_2_0_wb_clk_i),
    .Z(clknet_4_5_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_4_6_0_wb_clk_i (.I(clknet_3_3_0_wb_clk_i),
    .Z(clknet_4_6_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_4_7_0_wb_clk_i (.I(clknet_3_3_0_wb_clk_i),
    .Z(clknet_4_7_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_4_8_0_wb_clk_i (.I(clknet_3_4_0_wb_clk_i),
    .Z(clknet_4_8_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_4_9_0_wb_clk_i (.I(clknet_3_4_0_wb_clk_i),
    .Z(clknet_4_9_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_4_10_0_wb_clk_i (.I(clknet_3_5_0_wb_clk_i),
    .Z(clknet_4_10_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_4_11_0_wb_clk_i (.I(clknet_3_5_0_wb_clk_i),
    .Z(clknet_4_11_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_4_12_0_wb_clk_i (.I(clknet_3_6_0_wb_clk_i),
    .Z(clknet_4_12_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_4_13_0_wb_clk_i (.I(clknet_3_6_0_wb_clk_i),
    .Z(clknet_4_13_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_4_14_0_wb_clk_i (.I(clknet_3_7_0_wb_clk_i),
    .Z(clknet_4_14_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_4_15_0_wb_clk_i (.I(clknet_3_7_0_wb_clk_i),
    .Z(clknet_4_15_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_5_0_0_wb_clk_i (.I(clknet_4_0_0_wb_clk_i),
    .Z(clknet_5_0_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_5_1_0_wb_clk_i (.I(clknet_4_0_0_wb_clk_i),
    .Z(clknet_5_1_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_5_2_0_wb_clk_i (.I(clknet_4_1_0_wb_clk_i),
    .Z(clknet_5_2_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_5_3_0_wb_clk_i (.I(clknet_4_1_0_wb_clk_i),
    .Z(clknet_5_3_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_5_4_0_wb_clk_i (.I(clknet_4_2_0_wb_clk_i),
    .Z(clknet_5_4_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_5_5_0_wb_clk_i (.I(clknet_4_2_0_wb_clk_i),
    .Z(clknet_5_5_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_5_6_0_wb_clk_i (.I(clknet_4_3_0_wb_clk_i),
    .Z(clknet_5_6_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_5_7_0_wb_clk_i (.I(clknet_4_3_0_wb_clk_i),
    .Z(clknet_5_7_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_5_8_0_wb_clk_i (.I(clknet_4_4_0_wb_clk_i),
    .Z(clknet_5_8_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_5_9_0_wb_clk_i (.I(clknet_4_4_0_wb_clk_i),
    .Z(clknet_5_9_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_5_10_0_wb_clk_i (.I(clknet_4_5_0_wb_clk_i),
    .Z(clknet_5_10_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_5_11_0_wb_clk_i (.I(clknet_4_5_0_wb_clk_i),
    .Z(clknet_5_11_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_5_12_0_wb_clk_i (.I(clknet_4_6_0_wb_clk_i),
    .Z(clknet_5_12_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_5_13_0_wb_clk_i (.I(clknet_4_6_0_wb_clk_i),
    .Z(clknet_5_13_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_5_14_0_wb_clk_i (.I(clknet_4_7_0_wb_clk_i),
    .Z(clknet_5_14_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_5_15_0_wb_clk_i (.I(clknet_4_7_0_wb_clk_i),
    .Z(clknet_5_15_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_5_16_0_wb_clk_i (.I(clknet_4_8_0_wb_clk_i),
    .Z(clknet_5_16_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_5_17_0_wb_clk_i (.I(clknet_4_8_0_wb_clk_i),
    .Z(clknet_5_17_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_5_18_0_wb_clk_i (.I(clknet_4_9_0_wb_clk_i),
    .Z(clknet_5_18_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_5_19_0_wb_clk_i (.I(clknet_4_9_0_wb_clk_i),
    .Z(clknet_5_19_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_5_20_0_wb_clk_i (.I(clknet_4_10_0_wb_clk_i),
    .Z(clknet_5_20_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_5_21_0_wb_clk_i (.I(clknet_4_10_0_wb_clk_i),
    .Z(clknet_5_21_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_5_22_0_wb_clk_i (.I(clknet_4_11_0_wb_clk_i),
    .Z(clknet_5_22_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_5_23_0_wb_clk_i (.I(clknet_4_11_0_wb_clk_i),
    .Z(clknet_5_23_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_5_24_0_wb_clk_i (.I(clknet_4_12_0_wb_clk_i),
    .Z(clknet_5_24_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_5_25_0_wb_clk_i (.I(clknet_4_12_0_wb_clk_i),
    .Z(clknet_5_25_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_5_26_0_wb_clk_i (.I(clknet_4_13_0_wb_clk_i),
    .Z(clknet_5_26_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_5_27_0_wb_clk_i (.I(clknet_4_13_0_wb_clk_i),
    .Z(clknet_5_27_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_5_28_0_wb_clk_i (.I(clknet_4_14_0_wb_clk_i),
    .Z(clknet_5_28_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_5_29_0_wb_clk_i (.I(clknet_4_14_0_wb_clk_i),
    .Z(clknet_5_29_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_5_30_0_wb_clk_i (.I(clknet_4_15_0_wb_clk_i),
    .Z(clknet_5_30_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_5_31_0_wb_clk_i (.I(clknet_4_15_0_wb_clk_i),
    .Z(clknet_5_31_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_opt_1_0_wb_clk_i (.I(clknet_5_10_0_wb_clk_i),
    .Z(clknet_opt_1_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_opt_2_0_wb_clk_i (.I(clknet_5_11_0_wb_clk_i),
    .Z(clknet_opt_2_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_opt_3_0_wb_clk_i (.I(clknet_5_15_0_wb_clk_i),
    .Z(clknet_opt_3_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_opt_4_0_wb_clk_i (.I(clknet_5_15_0_wb_clk_i),
    .Z(clknet_opt_4_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_opt_5_0_wb_clk_i (.I(clknet_5_31_0_wb_clk_i),
    .Z(clknet_opt_5_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_1 (.I(_01551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_2 (.I(_02856_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_3 (.I(_02907_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_4 (.I(_05266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_5 (.I(\soc.rom_encoder_0.data_out[15] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_6 (.I(net15));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_7 (.I(net23));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_8 (.I(net28));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_9 (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_10 (.I(net76));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_11 (.I(net83));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_12 (.I(_02110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_13 (.I(\soc.cpu.AReg.data[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_14 (.I(net25));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_15 (.I(net44));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_16 (.I(net78));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1423 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1563 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1655 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1701 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_13 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_1_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_1_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_1_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_2_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_2_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_3_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_3_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_3_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_3_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_4_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_5_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_5_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_5_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_5_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_5_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_5_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_5_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_5_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_6_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_6_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_7_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_7_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_8_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_8_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_9_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_9_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_10_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_10_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_10_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_10_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_11_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_12_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_12_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_12_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_13_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_13_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_13_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_14_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_14_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_14_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_14_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_14_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_14_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_14_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_15_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_15_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_16_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_16_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_16_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_17_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_17_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_17_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_17_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_17_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_17_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_17_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_17_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_17_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_18_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_18_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_18_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_18_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_18_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_18_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_18_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_18_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_19_13 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_19_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_19_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_19_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_19_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_19_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_19_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_19_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_20_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_20_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_20_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_20_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_20_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_21_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_21_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_21_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_21_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_22_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_22_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_22_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_22_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_22_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_22_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_23_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_23_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_23_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_23_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_23_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1726 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_24_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_24_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_24_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_24_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_24_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_24_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_24_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_25_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_25_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_25_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_25_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_26_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_26_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_26_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_26_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_26_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_26_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_26_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_26_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_27_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_27_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_27_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_27_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_27_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_28_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_28_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_28_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_28_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_28_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_28_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_29_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_29_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_29_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_29_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_29_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_30_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_30_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_30_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_30_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_30_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_30_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_31_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_31_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_32_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_32_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_32_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_32_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_32_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1726 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_1743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_34_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_34_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_34_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_34_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_35_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_35_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_36_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_36_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_36_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_36_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_37_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_37_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_37_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_38_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_38_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_38_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_39_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_39_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_39_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_39_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_39_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_39_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_39_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_39_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_39_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_40_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_40_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_40_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_40_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_40_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_40_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_40_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_40_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_40_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_40_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_40_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_40_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_41_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_41_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_41_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_41_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_41_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_41_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_41_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_43_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_44_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_44_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_45_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_45_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_45_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_45_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_45_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_45_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_46_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_47_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_1384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_47_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_47_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_48_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_48_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_1702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_49_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_49_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_49_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_50_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_50_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_51_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_51_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_52_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_52_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_52_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1423 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_1440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_1508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_53_1385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1726 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_54_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_54_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_1440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_55_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_55_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_56_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_56_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_57_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_57_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_58_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_58_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_58_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_1702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_59_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_59_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_60_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_60_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_60_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1423 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_60_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_60_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_1702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_61_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_1458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_61_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_62_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_62_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_1514 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_63_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_1481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_63_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_64_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_64_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_65_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_1532 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_1548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_65_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_66_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_66_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_66_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_67_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_1483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_1513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_1545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_67_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_68_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_69_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_69_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_1509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_69_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_70_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_71_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_1534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_1550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_71_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_72_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_72_1535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_1583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_1509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_73_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_73_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_74_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_74_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_75_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_75_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_1483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_75_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_76_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_77_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_77_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_78_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1421 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_79_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_1474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_1533 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_1549 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_79_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_80_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_80_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_80_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_1518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_80_1535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_1583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_81_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_81_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_81_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_81_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_82_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1423 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_82_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_83_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_83_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1462 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_1548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_83_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_84_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_84_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_84_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_84_1535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_1583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_85_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_85_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_85_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_85_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_86_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_86_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_86_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1532 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_86_1548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_87_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_87_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_1478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_87_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_88_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_88_1474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_1506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_88_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_89_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_89_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1455 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_1509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_1546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_89_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_90_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_90_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_90_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_1702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_91_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_91_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_91_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1532 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_92_1549 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_93_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_1615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1631 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_93_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_94_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_1435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_1508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_94_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_1589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_1543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_95_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_96_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1532 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_96_1563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_97_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_1526 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_1549 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_97_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_98_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_98_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_98_1479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_1517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_99_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_1535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_1551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_99_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_100_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_100_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1423 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_1518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_100_1535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_1583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_101_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_1471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_1545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_101_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_103_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_1543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_103_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_104_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_1518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_104_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_105_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_105_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_106_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1532 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_106_1548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_1483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_107_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_108_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_108_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_108_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_109_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_109_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_109_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_1483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_109_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1726 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_1743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_110_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_1440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_1509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_111_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1385 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_111_1517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_1549 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_111_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_112_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_1515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_112_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_112_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_1702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_113_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1458 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1526 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_113_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_114_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_114_1478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_1510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_114_1535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_1583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_115_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_116_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_116_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_1505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_117_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_118_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_118_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_118_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_118_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_118_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_119_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_119_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_1462 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_1478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_119_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_120_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_120_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_120_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_120_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_120_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_120_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_1508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_121_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_121_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_122_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_123_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_1483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_123_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_124_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_124_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_1505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_126_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_126_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_127_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_127_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_127_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_128_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_129_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_129_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_129_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_129_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_131_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_131_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_132_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_132_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_132_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_132_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_132_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_1702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_133_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_134_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_134_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_134_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_135_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_135_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_135_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_136_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_136_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_136_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_136_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_136_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_136_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_137_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_137_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_137_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_137_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_137_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_137_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_137_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_137_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_137_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_138_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_138_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_138_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_138_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_138_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_138_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_138_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_139_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_139_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_139_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_139_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_139_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_139_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_139_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_139_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_139_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_140_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_140_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_140_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_140_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_141_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_141_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_141_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_141_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_141_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_141_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_141_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_141_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_141_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_141_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_141_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_141_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_142_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_142_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_142_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_142_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_142_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_143_13 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_143_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_143_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_143_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_144_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_145_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_145_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_145_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_145_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_145_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_145_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_145_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_145_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_145_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_145_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_145_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_145_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_145_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_145_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_145_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_145_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_145_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_145_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_145_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_145_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_146_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_146_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_146_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_146_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_146_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_146_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_146_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_146_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_146_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_146_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_146_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_146_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_146_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_146_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_146_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_146_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_1753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_146_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_147_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_147_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_147_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_147_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_147_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_147_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_147_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_147_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_147_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_147_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_147_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_147_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_147_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_147_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_147_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_147_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_147_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_147_1722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_147_1726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_1728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_147_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_148_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_148_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_148_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_148_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_148_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_148_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_148_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_148_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_148_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_148_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_148_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_148_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_148_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_148_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_148_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_148_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_1420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_1423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_148_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_148_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_148_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_148_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_148_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_149_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_149_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_149_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_149_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_149_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_149_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_149_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_149_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_149_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_149_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_149_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_149_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_149_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_149_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_149_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_149_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_149_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_149_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_149_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_149_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_149_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_150_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_150_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_150_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_150_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_150_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_150_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_150_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_150_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_150_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_150_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_150_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_150_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_150_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_150_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_150_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_150_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_150_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_150_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_150_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_150_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_150_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_150_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_150_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_150_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_150_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_151_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_151_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_151_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_151_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_151_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_151_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_151_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_151_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_151_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_151_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_151_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_151_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_151_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_151_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_151_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_151_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_151_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_151_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_152_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_152_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_152_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_152_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_152_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_152_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_152_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_152_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_152_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_152_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_152_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_152_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_152_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_152_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_152_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_152_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_152_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_152_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_152_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_152_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_152_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_153_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_153_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_153_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_153_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_153_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_153_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_153_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_153_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_153_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_153_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_153_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_153_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_153_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_153_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_153_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_153_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_153_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_153_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_153_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_1384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_153_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_153_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_153_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_153_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_153_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_154_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_154_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_154_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_154_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_154_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_154_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_154_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_154_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_154_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_154_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_154_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_154_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_154_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_154_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_154_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_154_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_154_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_154_1702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_154_1718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_154_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_154_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_154_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_155_13 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_155_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_155_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_155_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_155_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_155_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_155_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_155_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_155_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_155_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_155_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_155_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_155_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_155_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_155_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_155_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_155_1462 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_155_1478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_155_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_155_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_155_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_155_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_155_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_156_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_156_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_156_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_156_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_156_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_156_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_156_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_156_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_156_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_156_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_156_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_156_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_156_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_156_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_156_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_156_1678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_1680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_156_1731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_156_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_156_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_1753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_156_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_157_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_157_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_157_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_157_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_157_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_157_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_157_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_157_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_157_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_157_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_157_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_157_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_157_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_157_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_157_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_157_1722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_157_1726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_1728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_157_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_158_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_158_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_158_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_158_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_158_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_158_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_158_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_158_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_158_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_158_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_158_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_158_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_158_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_158_1435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_158_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_158_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_158_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_158_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_158_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_159_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_159_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_159_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_159_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_159_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_159_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_159_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_159_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_159_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_159_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_159_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_159_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_159_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_159_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_159_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_159_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_159_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_160_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_160_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_160_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_160_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_160_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_160_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_160_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_160_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_160_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_160_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_160_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_160_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_160_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_160_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_160_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_161_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_161_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_161_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_161_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_161_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_161_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_161_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_161_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_161_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_161_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_161_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_161_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_161_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_162_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_162_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_162_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_162_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_162_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_162_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_162_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_162_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_162_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_162_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_162_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_162_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_162_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_162_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_162_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_162_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_162_1702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_162_1718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_1722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_162_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_162_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_162_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_163_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_163_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_163_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_163_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_163_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_163_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_163_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_163_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_163_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_163_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_163_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_163_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_163_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_163_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_163_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_164_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_164_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_164_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_164_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_164_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_164_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_164_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_164_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_164_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_164_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_165_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_165_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_165_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_165_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_165_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_165_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_165_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_165_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_165_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_165_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_165_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_165_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_165_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_166_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_166_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_166_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_166_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_166_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_166_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_166_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_166_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_166_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_166_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_166_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_166_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_166_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_166_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_166_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_166_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_166_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_166_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_166_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_166_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_166_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_167_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_167_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_167_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_167_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_167_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_167_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_167_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_167_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_167_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_167_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_167_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_167_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_167_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_167_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_167_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_167_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_168_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_168_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_168_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_168_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_168_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_168_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_168_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_168_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_168_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_168_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_168_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_168_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_168_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_168_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_168_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_169_13 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_169_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_169_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_169_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_169_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_169_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_169_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_169_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_169_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_169_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_169_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_169_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_169_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_169_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_169_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_169_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_169_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_169_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_169_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_169_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_169_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_170_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_170_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_170_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_170_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_170_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_170_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_170_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_170_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_170_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_170_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_170_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_170_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_170_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_170_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_170_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_170_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_170_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_170_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_170_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_170_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_170_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_170_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_170_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_171_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_171_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_171_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_171_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_171_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_171_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_171_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_171_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_171_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_171_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_171_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_171_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_171_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_171_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_171_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_171_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_171_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_171_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_171_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_171_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_171_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_172_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_172_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_172_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_172_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_172_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_172_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_172_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_172_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_172_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_172_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_172_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_172_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_172_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_172_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_172_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_172_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_172_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_172_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_172_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_172_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_173_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_173_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_173_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_173_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_173_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_173_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_173_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_173_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_173_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_173_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_173_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_173_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_173_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_173_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_173_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_173_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_173_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_173_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_173_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_173_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_174_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_174_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_174_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_174_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_174_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_174_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_174_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_174_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_174_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_174_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_174_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_174_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_174_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_174_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_174_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_174_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_1753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_174_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_175_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_175_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_175_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_175_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_175_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_175_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_175_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_175_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_175_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_175_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_175_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_175_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_175_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_175_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_175_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_175_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_175_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_175_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_175_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_175_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_175_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_176_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_176_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_176_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_176_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_176_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_176_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_176_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_176_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_176_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_176_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_176_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_176_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_176_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_176_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_176_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_176_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_176_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_176_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_176_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_176_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_176_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_176_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_176_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_1448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_176_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_176_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_176_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_176_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_176_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_176_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_176_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_1753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_176_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_177_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_177_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_177_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_177_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_177_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_177_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_177_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_177_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_177_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_177_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_177_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_177_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_177_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_177_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_177_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_177_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_178_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_178_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_178_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_178_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_178_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_178_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_178_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_178_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_178_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_178_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_178_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_178_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_178_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_178_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_178_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_178_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_179_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_179_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_179_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_179_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_179_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_179_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_179_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_179_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_179_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_179_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_180_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_180_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_180_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_180_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_180_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_180_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_180_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_180_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_180_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_180_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_180_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_180_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_180_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_180_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_180_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_180_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_180_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_180_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_180_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_180_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_181_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_181_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_181_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_181_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_181_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_181_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_181_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_181_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_181_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_181_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_181_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_181_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_181_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_181_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_181_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_182_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_182_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_182_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_182_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_182_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_182_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_182_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_182_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_182_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_182_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_182_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_182_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_182_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_182_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_182_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_182_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_183_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_183_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_183_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_183_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_183_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_183_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_183_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_183_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_183_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_183_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_183_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_183_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_183_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_183_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_183_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_183_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_183_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_183_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_183_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_184_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_184_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_184_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_184_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_184_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_184_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_184_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_184_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_184_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_184_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_184_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_184_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_184_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_184_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_184_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_184_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_184_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_184_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_184_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_184_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_184_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_184_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_184_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_184_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_184_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_184_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_184_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_184_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_184_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_184_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_184_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_184_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_184_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_184_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_184_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_184_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_185_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_185_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_185_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_185_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_185_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_185_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_185_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_185_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_185_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_185_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_185_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_185_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_185_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_185_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_185_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_185_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_185_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_185_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_185_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_185_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_185_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_185_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_185_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_185_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_185_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_185_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_185_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_185_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_185_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_185_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_185_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_185_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_185_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_185_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_185_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_185_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_185_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_185_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_185_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_185_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_186_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_186_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_186_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_186_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_186_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_186_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_186_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_186_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_186_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_186_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_186_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_186_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_186_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_186_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_186_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_186_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_186_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_186_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_186_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_186_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_186_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_186_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_186_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_186_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_186_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_186_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_186_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_186_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_186_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_186_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_186_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_186_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_186_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_186_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_186_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_186_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_186_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_186_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_186_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_1753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_186_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_187_13 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_187_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_187_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_187_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_187_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_187_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_187_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_187_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_187_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_187_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_187_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_187_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_187_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_187_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_187_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_187_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_187_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_187_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_187_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_187_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_187_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_187_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_187_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_187_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_187_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_187_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_187_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_187_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_187_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_187_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_187_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_187_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_187_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_187_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_187_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_188_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_188_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_188_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_188_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_188_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_188_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_188_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_188_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_188_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_188_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_188_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_188_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_188_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_188_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_188_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_188_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_188_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_188_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_188_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_188_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_188_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_188_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_188_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_188_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_188_1702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_188_1718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_188_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_188_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_188_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_189_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_189_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_189_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_189_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_189_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_189_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_189_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_189_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_189_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_189_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_189_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_189_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_189_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_189_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_189_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_189_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_189_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_189_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_190_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_190_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_190_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_190_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_190_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_190_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_190_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_190_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_190_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_190_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_190_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_190_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_190_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_190_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_190_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_190_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_190_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_190_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_190_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_190_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_191_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_191_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_191_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_191_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_191_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_191_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_191_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_191_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_191_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_191_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_191_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_191_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_191_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_191_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_191_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_191_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_191_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_191_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_191_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_192_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_192_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_192_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_192_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_192_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_192_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_192_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_192_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_192_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_192_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_192_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_192_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_192_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_192_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_192_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_193_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_193_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_193_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_193_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_193_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_193_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_193_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_193_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_193_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_193_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_193_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_193_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_193_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_193_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_194_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_194_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_194_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_194_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_194_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_194_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_194_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_194_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_194_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_194_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_194_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_194_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_194_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_194_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_195_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_195_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_195_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_195_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_195_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_195_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_195_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_195_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_195_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_195_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_195_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_195_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_195_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_195_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_195_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_195_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_195_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_195_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_195_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_195_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_195_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_195_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_195_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_195_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_195_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_195_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_195_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_195_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_196_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_196_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_196_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_196_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_196_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_196_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_196_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_196_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_196_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_196_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_196_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_196_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_196_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_196_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_196_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_196_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_196_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_196_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_196_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_196_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_196_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_196_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_196_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_196_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_196_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_196_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_196_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_196_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_196_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_197_13 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_197_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_197_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_197_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_197_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_197_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_197_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_197_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_197_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_197_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_197_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_197_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_197_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_197_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_197_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_197_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_197_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_197_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_197_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_197_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_197_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_197_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_197_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_197_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_197_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_197_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_197_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_197_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_197_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_197_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_197_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_198_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_198_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_198_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_198_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_198_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_198_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_198_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_198_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_198_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_198_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_198_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_198_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_198_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_198_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_198_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_198_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_198_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_198_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_198_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_198_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_198_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_198_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_198_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_198_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_198_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_198_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_198_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_198_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_1753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_198_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_199_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_199_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_199_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_199_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_199_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_199_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_199_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_199_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_199_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_199_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_199_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_199_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_199_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_199_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_199_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_199_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_199_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_199_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_199_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_199_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_199_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_199_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_199_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_199_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_199_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_199_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_199_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_199_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_200_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_200_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_200_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_200_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_200_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_200_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_200_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_200_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_200_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_200_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_200_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_200_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_200_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_200_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_200_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_200_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_200_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_200_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_200_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_200_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_200_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_200_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_200_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_200_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_200_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_200_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_200_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_200_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_200_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_201_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_201_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_201_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_201_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_201_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_201_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_201_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_201_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_201_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_201_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_201_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_201_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_201_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_201_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_201_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_201_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_201_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_201_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_201_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_201_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_201_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_201_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_201_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_201_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_201_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_201_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_201_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_201_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_202_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_202_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_202_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_202_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_202_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_202_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_202_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_202_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_202_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_202_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_202_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_202_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_202_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_202_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_202_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_202_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_202_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_202_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_202_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_202_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_202_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_202_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_202_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_202_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_202_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_202_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_202_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_202_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_202_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_203_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_203_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_203_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_203_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_203_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_203_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_203_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_203_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_203_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_203_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_203_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_203_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_203_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_203_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_203_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_203_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_203_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_203_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_203_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_203_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_203_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_203_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_203_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_203_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_203_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_203_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_203_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_203_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_204_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_204_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_204_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_204_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_204_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_204_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_204_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_204_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_204_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_204_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_204_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_204_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_204_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_204_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_204_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_204_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_204_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_204_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_204_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_204_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_204_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_204_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_204_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_204_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_204_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_204_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_204_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_204_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_204_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_205_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_205_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_205_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_205_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_205_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_205_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_205_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_205_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_205_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_205_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_205_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_205_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_205_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_205_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_205_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_205_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_205_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_205_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_205_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_205_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_205_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_205_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_205_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_205_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_205_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_205_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_205_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_205_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_206_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_206_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_206_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_206_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_206_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_206_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_206_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_206_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_206_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_206_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_206_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_206_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_206_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_206_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_206_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_206_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_206_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_206_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_206_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_206_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_206_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_206_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_206_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_206_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_206_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_206_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_206_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_206_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_206_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_207_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_207_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_207_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_207_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_207_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_207_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_207_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_207_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_207_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_207_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_207_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_207_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_207_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_207_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_207_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_207_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_207_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_207_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_207_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_207_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_207_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_207_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_207_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_207_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_207_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_207_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_207_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_207_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_208_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_208_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_208_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_208_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_208_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_208_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_208_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_208_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_208_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_208_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_208_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_208_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_208_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_208_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_208_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_208_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_208_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_208_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_208_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_208_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_208_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_208_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_208_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_208_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_208_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_208_1702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_208_1718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_208_1722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_208_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_208_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_208_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_209_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_209_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_209_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_209_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_209_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_209_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_209_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_209_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_209_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_209_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_209_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_209_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_209_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_209_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_209_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_209_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_209_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_209_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_209_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_209_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_209_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_209_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_209_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_209_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_209_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_209_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_209_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_209_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_210_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_210_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_210_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_210_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_210_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_210_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_210_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_210_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_210_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_210_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_210_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_210_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_210_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_210_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_210_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_210_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_210_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_210_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_210_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_210_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_210_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_210_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_210_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_210_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_210_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_210_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_210_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_210_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_1753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_210_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_211_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_211_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_211_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_211_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_211_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_211_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_211_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_211_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_211_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_211_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_211_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_211_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_211_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_211_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_211_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_211_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_211_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_211_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_211_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_211_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_211_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_211_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_211_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_211_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_211_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_211_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_211_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_211_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_212_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_212_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_212_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_212_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_212_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_212_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_212_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_212_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_212_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_212_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_212_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_212_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_212_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_212_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_212_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_212_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_212_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_212_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_212_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_212_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_212_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_212_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_212_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_212_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_212_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_212_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_212_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_212_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_212_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_213_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_213_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_213_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_213_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_213_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_213_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_213_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_213_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_213_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_213_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_213_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_213_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_213_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_213_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_213_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_213_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_213_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_213_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_213_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_213_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_213_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_213_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_213_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_213_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_213_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_213_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_213_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_213_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_214_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_214_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_214_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_214_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_214_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_214_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_214_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_214_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_214_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_214_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_214_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_214_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_214_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_214_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_214_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_214_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_214_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_214_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_214_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_214_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_214_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_214_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_214_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_214_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_214_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_214_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_214_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_214_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_214_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_215_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_215_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_215_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_215_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_215_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_215_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_215_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_215_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_215_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_215_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_215_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_215_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_215_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_215_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_215_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_215_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_215_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_215_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_215_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_215_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_215_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_215_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_215_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_215_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_215_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_215_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_215_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_215_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_216_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_216_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_216_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_216_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_216_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_216_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_216_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_216_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_216_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_216_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_216_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_216_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_216_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_216_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_216_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_216_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_216_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_216_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_216_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_216_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_216_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_216_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_216_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_216_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_216_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_216_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_216_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_216_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_216_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_217_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_217_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_217_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_217_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_217_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_217_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_217_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_217_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_217_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_217_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_217_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_217_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_217_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_217_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_217_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_217_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_217_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_217_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_217_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_217_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_217_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_217_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_217_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_217_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_217_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_217_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_217_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_217_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_218_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_218_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_218_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_218_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_218_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_218_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_218_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_218_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_218_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_218_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_218_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_218_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_218_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_218_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_218_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_218_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_218_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_218_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_218_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_218_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_218_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_218_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_218_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_218_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_218_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_218_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_218_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_218_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_218_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_219_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_219_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_219_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_219_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_219_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_219_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_219_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_219_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_219_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_219_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_219_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_219_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_219_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_219_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_219_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_219_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_219_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_219_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_219_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_219_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_219_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_219_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_219_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_219_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_219_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_219_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_219_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_219_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_220_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_220_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_220_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_220_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_220_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_220_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_220_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_220_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_220_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_220_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_220_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_220_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_220_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_220_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_220_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_220_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_220_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_220_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_220_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_220_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_220_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_220_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_220_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_220_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_220_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_220_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_220_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_220_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_220_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_221_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_221_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_221_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_221_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_221_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_221_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_221_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_221_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_221_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_221_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_221_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_221_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_221_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_221_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_221_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_221_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_221_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_221_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_221_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_221_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_221_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_221_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_221_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_221_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_221_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_221_1722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_221_1726 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_221_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_221_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_222_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_222_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_222_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_222_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_222_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_222_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_222_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_222_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_222_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_222_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_222_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_222_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_222_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_222_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_222_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_222_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_222_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_222_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_222_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_222_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_222_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_222_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_222_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_222_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_222_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_222_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_222_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_1753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_222_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_223_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_223_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_223_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_223_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_223_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_223_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_223_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_223_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_223_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_223_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_223_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_223_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_223_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_223_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_223_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_223_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_223_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_223_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_223_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_223_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_223_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_223_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_223_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_223_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_223_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_223_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_223_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_223_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_224_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_224_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_224_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_224_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_224_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_224_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_224_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_224_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_224_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_224_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_224_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_224_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_224_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_224_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_224_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_224_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_224_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_224_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_224_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_224_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_224_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_224_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_224_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_224_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_224_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_224_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_224_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_224_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_224_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_225_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_225_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_225_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_225_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_225_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_225_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_225_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_225_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_225_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_225_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_225_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_225_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_225_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_225_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_225_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_225_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_225_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_225_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_225_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_225_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_225_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_225_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_225_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_225_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_225_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_225_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_225_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_225_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_226_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_226_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_226_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_226_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_226_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_226_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_226_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_226_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_226_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_226_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_226_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_226_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_226_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_226_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_226_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_226_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_226_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_226_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_226_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_226_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_226_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_226_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_226_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_226_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_226_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_226_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_226_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_226_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_226_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_227_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_227_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_227_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_227_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_227_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_227_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_227_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_227_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_227_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_227_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_227_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_227_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_227_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_227_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_227_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_227_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_227_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_227_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_227_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_227_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_227_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_227_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_227_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_227_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_227_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_227_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_227_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_227_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_227_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_228_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_228_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_228_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_228_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_228_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_228_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_228_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_228_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_228_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_228_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_228_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_228_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_228_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_228_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_228_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_228_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_228_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_228_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_228_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_228_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_228_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_228_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_228_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_228_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_228_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_228_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_228_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_228_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_228_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_229_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_229_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_229_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_229_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_229_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_229_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_229_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_229_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_229_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_229_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_229_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_229_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_229_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_229_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_229_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_229_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_229_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_229_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_229_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_229_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_229_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_229_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_229_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_229_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_229_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_229_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_229_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_229_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_230_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_230_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_230_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_230_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_230_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_230_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_230_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_230_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_230_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_230_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_230_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_230_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_230_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_230_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_230_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_230_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_230_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_230_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_230_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_230_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_230_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_230_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_230_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_230_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_230_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_230_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_230_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_1753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_230_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_231_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_231_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_231_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_231_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_231_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_231_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_231_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_231_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_231_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_231_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_231_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_231_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_231_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_231_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_231_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_231_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_231_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_231_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_231_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_231_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_231_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_231_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_231_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_231_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_231_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_231_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_231_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_231_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_232_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_232_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_232_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_232_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_232_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_232_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_232_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_232_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_232_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_232_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_232_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_232_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_232_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_232_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_232_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_232_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_232_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_232_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_232_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_232_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_232_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_232_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_232_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_232_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_232_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_232_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_232_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_232_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_232_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_233_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_233_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_233_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_233_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_233_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_233_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_233_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_233_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_233_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_233_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_233_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_233_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_233_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_233_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_233_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_233_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_233_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_233_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_233_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_233_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_233_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_233_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_233_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_233_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_233_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_233_1722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_233_1726 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_233_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_233_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_234_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_234_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_234_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_234_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_234_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_234_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_234_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_234_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_234_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_234_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_234_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_234_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_234_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_234_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_234_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_234_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_234_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_234_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_234_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_234_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_234_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_234_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_234_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_234_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_234_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_234_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_234_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_234_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_234_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_234_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_235_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_235_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_235_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_235_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_235_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_235_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_235_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_235_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_235_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_235_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_235_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_235_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_235_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_235_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_235_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_235_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_235_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_235_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_235_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_235_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_235_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_235_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_235_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_235_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_235_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_235_1722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_235_1726 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_235_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_235_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_236_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_236_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_236_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_236_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_236_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_236_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_236_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_236_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_236_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_236_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_236_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_236_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_236_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_236_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_236_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_236_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_236_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_236_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_236_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_236_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_236_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_236_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_236_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_236_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_236_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_236_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_236_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_236_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_236_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_237_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_237_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_237_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_237_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_237_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_237_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_237_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_237_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_237_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_237_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_237_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_237_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_237_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_237_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_237_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_237_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_237_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_237_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_237_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_237_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_237_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_237_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_237_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_237_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_237_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_237_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_237_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_237_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_238_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_238_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_238_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_238_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_238_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_238_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_238_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_238_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_238_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_238_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_238_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_238_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_238_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_238_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_238_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_238_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_238_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_238_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_238_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_238_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_238_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_238_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_238_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_238_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_238_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_238_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_238_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_238_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_238_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_239_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_239_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_239_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_239_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_239_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_239_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_239_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_239_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_239_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_239_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_239_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_239_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_239_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_239_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_239_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_239_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_239_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_239_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_239_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_239_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_239_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_239_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_239_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_239_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_239_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_239_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_239_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_239_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_240_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_240_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_240_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_240_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_240_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_240_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_240_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_240_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_240_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_240_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_240_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_240_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_240_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_240_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_240_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_240_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_240_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_240_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_240_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_240_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_240_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_240_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_240_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_240_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_240_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_240_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_240_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_240_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_240_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_241_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_241_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_241_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_241_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_241_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_241_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_241_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_241_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_241_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_241_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_241_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_241_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_241_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_241_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_241_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_241_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_241_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_241_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_241_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_241_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_241_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_241_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_241_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_241_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_241_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_241_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_241_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_241_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_242_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_242_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_242_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_242_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_242_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_242_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_242_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_242_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_242_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_242_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_242_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_242_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_242_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_242_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_242_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_242_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_242_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_242_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_242_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_242_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_242_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_242_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_242_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_242_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_242_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_242_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_242_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_242_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_1753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_242_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_243_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_243_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_243_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_243_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_243_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_243_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_243_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_243_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_243_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_243_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_243_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_243_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_243_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_243_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_243_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_243_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_243_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_243_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_243_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_243_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_243_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_243_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_243_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_243_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_243_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_243_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_243_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_243_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_244_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_244_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_244_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_244_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_244_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_244_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_244_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_244_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_244_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_244_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_244_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_244_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_244_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_244_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_244_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_244_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_244_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_244_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_244_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_244_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_244_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_244_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_244_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_244_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_244_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_244_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_244_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_244_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_244_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_244_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_244_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_245_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_245_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_245_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_245_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_245_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_245_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_245_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_245_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_245_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_245_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_245_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_245_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_245_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_245_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_245_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_245_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_245_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_245_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_245_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_245_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_245_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_245_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_245_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_245_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_245_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_245_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_245_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_245_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_245_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_1442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_245_1448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_245_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_245_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_245_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_245_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_245_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_245_1722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_245_1726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_245_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_13 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_246_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_246_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_246_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_246_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_246_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_246_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_246_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_246_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_246_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_246_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_246_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_246_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_246_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_246_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_246_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_246_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_246_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_246_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_246_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_246_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_246_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_246_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_246_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_246_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_246_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_246_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_246_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_246_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_246_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_246_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_246_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_246_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_246_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_246_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_246_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_246_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_246_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_246_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_246_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_246_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_246_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_246_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_246_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_246_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_246_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_246_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_246_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_246_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_246_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_246_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_246_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_246_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_246_1442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_246_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_246_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_246_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_246_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_246_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_246_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_1620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_1624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_1626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_246_1631 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_246_1639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_1643 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_246_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_246_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_1714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_246_1742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_246_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_246_1757 ();
 assign io_oeb[0] = net91;
 assign io_oeb[14] = net101;
 assign io_oeb[15] = net102;
 assign io_oeb[1] = net92;
 assign io_oeb[20] = net103;
 assign io_oeb[21] = net104;
 assign io_oeb[26] = net224;
 assign io_oeb[27] = net105;
 assign io_oeb[28] = net106;
 assign io_oeb[29] = net107;
 assign io_oeb[2] = net93;
 assign io_oeb[30] = net225;
 assign io_oeb[31] = net226;
 assign io_oeb[32] = net227;
 assign io_oeb[33] = net228;
 assign io_oeb[34] = net108;
 assign io_oeb[35] = net109;
 assign io_oeb[36] = net110;
 assign io_oeb[37] = net111;
 assign io_oeb[3] = net94;
 assign io_oeb[4] = net95;
 assign io_oeb[5] = net96;
 assign io_oeb[6] = net97;
 assign io_oeb[7] = net98;
 assign io_oeb[8] = net99;
 assign io_oeb[9] = net100;
 assign io_out[0] = net112;
 assign io_out[1] = net113;
 assign io_out[26] = net120;
 assign io_out[2] = net114;
 assign io_out[30] = net121;
 assign io_out[31] = net122;
 assign io_out[32] = net123;
 assign io_out[33] = net124;
 assign io_out[3] = net115;
 assign io_out[4] = net116;
 assign io_out[5] = net117;
 assign io_out[6] = net118;
 assign io_out[7] = net119;
 assign irq[0] = net125;
 assign irq[1] = net126;
 assign irq[2] = net127;
 assign la_data_out[0] = net128;
 assign la_data_out[10] = net138;
 assign la_data_out[11] = net139;
 assign la_data_out[12] = net140;
 assign la_data_out[13] = net141;
 assign la_data_out[14] = net142;
 assign la_data_out[15] = net143;
 assign la_data_out[16] = net144;
 assign la_data_out[17] = net145;
 assign la_data_out[18] = net146;
 assign la_data_out[19] = net147;
 assign la_data_out[1] = net129;
 assign la_data_out[20] = net148;
 assign la_data_out[21] = net149;
 assign la_data_out[22] = net150;
 assign la_data_out[23] = net151;
 assign la_data_out[24] = net152;
 assign la_data_out[25] = net153;
 assign la_data_out[26] = net154;
 assign la_data_out[28] = net155;
 assign la_data_out[29] = net156;
 assign la_data_out[2] = net130;
 assign la_data_out[30] = net157;
 assign la_data_out[31] = net158;
 assign la_data_out[32] = net159;
 assign la_data_out[33] = net160;
 assign la_data_out[34] = net161;
 assign la_data_out[35] = net162;
 assign la_data_out[36] = net163;
 assign la_data_out[37] = net164;
 assign la_data_out[38] = net165;
 assign la_data_out[39] = net166;
 assign la_data_out[3] = net131;
 assign la_data_out[40] = net167;
 assign la_data_out[41] = net168;
 assign la_data_out[42] = net169;
 assign la_data_out[43] = net170;
 assign la_data_out[44] = net171;
 assign la_data_out[45] = net172;
 assign la_data_out[46] = net173;
 assign la_data_out[47] = net174;
 assign la_data_out[48] = net175;
 assign la_data_out[49] = net176;
 assign la_data_out[4] = net132;
 assign la_data_out[50] = net177;
 assign la_data_out[51] = net178;
 assign la_data_out[52] = net179;
 assign la_data_out[53] = net180;
 assign la_data_out[54] = net181;
 assign la_data_out[55] = net182;
 assign la_data_out[56] = net183;
 assign la_data_out[57] = net184;
 assign la_data_out[58] = net185;
 assign la_data_out[59] = net186;
 assign la_data_out[5] = net133;
 assign la_data_out[60] = net187;
 assign la_data_out[61] = net188;
 assign la_data_out[62] = net189;
 assign la_data_out[63] = net190;
 assign la_data_out[6] = net134;
 assign la_data_out[7] = net135;
 assign la_data_out[8] = net136;
 assign la_data_out[9] = net137;
 assign wbs_ack_o = net191;
 assign wbs_dat_o[0] = net192;
 assign wbs_dat_o[10] = net202;
 assign wbs_dat_o[11] = net203;
 assign wbs_dat_o[12] = net204;
 assign wbs_dat_o[13] = net205;
 assign wbs_dat_o[14] = net206;
 assign wbs_dat_o[15] = net207;
 assign wbs_dat_o[16] = net208;
 assign wbs_dat_o[17] = net209;
 assign wbs_dat_o[18] = net210;
 assign wbs_dat_o[19] = net211;
 assign wbs_dat_o[1] = net193;
 assign wbs_dat_o[20] = net212;
 assign wbs_dat_o[21] = net213;
 assign wbs_dat_o[22] = net214;
 assign wbs_dat_o[23] = net215;
 assign wbs_dat_o[24] = net216;
 assign wbs_dat_o[25] = net217;
 assign wbs_dat_o[26] = net218;
 assign wbs_dat_o[27] = net219;
 assign wbs_dat_o[28] = net220;
 assign wbs_dat_o[29] = net221;
 assign wbs_dat_o[2] = net194;
 assign wbs_dat_o[30] = net222;
 assign wbs_dat_o[31] = net223;
 assign wbs_dat_o[3] = net195;
 assign wbs_dat_o[4] = net196;
 assign wbs_dat_o[5] = net197;
 assign wbs_dat_o[6] = net198;
 assign wbs_dat_o[7] = net199;
 assign wbs_dat_o[8] = net200;
 assign wbs_dat_o[9] = net201;
endmodule

