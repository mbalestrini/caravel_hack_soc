// This is the unpowered netlist.
module caravel_hack_soc (wb_clk_i,
    wb_rst_i,
    wbs_ack_o,
    wbs_cyc_i,
    wbs_stb_i,
    wbs_we_i,
    io_in,
    io_oeb,
    io_out,
    irq,
    la_data_in,
    la_data_out,
    la_oenb,
    wbs_adr_i,
    wbs_dat_i,
    wbs_dat_o,
    wbs_sel_i);
 input wb_clk_i;
 input wb_rst_i;
 output wbs_ack_o;
 input wbs_cyc_i;
 input wbs_stb_i;
 input wbs_we_i;
 input [37:0] io_in;
 output [37:0] io_oeb;
 output [37:0] io_out;
 output [2:0] irq;
 input [63:0] la_data_in;
 output [63:0] la_data_out;
 input [63:0] la_oenb;
 input [31:0] wbs_adr_i;
 input [31:0] wbs_dat_i;
 output [31:0] wbs_dat_o;
 input [3:0] wbs_sel_i;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire _2063_;
 wire _2064_;
 wire _2065_;
 wire _2066_;
 wire _2067_;
 wire _2068_;
 wire _2069_;
 wire _2070_;
 wire _2071_;
 wire _2072_;
 wire _2073_;
 wire _2074_;
 wire _2075_;
 wire _2076_;
 wire _2077_;
 wire _2078_;
 wire _2079_;
 wire _2080_;
 wire _2081_;
 wire _2082_;
 wire _2083_;
 wire _2084_;
 wire _2085_;
 wire _2086_;
 wire _2087_;
 wire _2088_;
 wire _2089_;
 wire _2090_;
 wire _2091_;
 wire _2092_;
 wire _2093_;
 wire _2094_;
 wire _2095_;
 wire _2096_;
 wire _2097_;
 wire _2098_;
 wire _2099_;
 wire _2100_;
 wire _2101_;
 wire _2102_;
 wire _2103_;
 wire _2104_;
 wire _2105_;
 wire _2106_;
 wire _2107_;
 wire _2108_;
 wire _2109_;
 wire _2110_;
 wire _2111_;
 wire _2112_;
 wire _2113_;
 wire _2114_;
 wire _2115_;
 wire _2116_;
 wire _2117_;
 wire _2118_;
 wire _2119_;
 wire _2120_;
 wire _2121_;
 wire _2122_;
 wire _2123_;
 wire _2124_;
 wire _2125_;
 wire _2126_;
 wire _2127_;
 wire _2128_;
 wire _2129_;
 wire _2130_;
 wire _2131_;
 wire _2132_;
 wire _2133_;
 wire _2134_;
 wire _2135_;
 wire _2136_;
 wire _2137_;
 wire _2138_;
 wire _2139_;
 wire _2140_;
 wire _2141_;
 wire _2142_;
 wire _2143_;
 wire _2144_;
 wire _2145_;
 wire _2146_;
 wire _2147_;
 wire _2148_;
 wire _2149_;
 wire _2150_;
 wire _2151_;
 wire _2152_;
 wire _2153_;
 wire _2154_;
 wire _2155_;
 wire _2156_;
 wire _2157_;
 wire _2158_;
 wire _2159_;
 wire _2160_;
 wire _2161_;
 wire _2162_;
 wire _2163_;
 wire _2164_;
 wire _2165_;
 wire _2166_;
 wire _2167_;
 wire _2168_;
 wire _2169_;
 wire _2170_;
 wire _2171_;
 wire _2172_;
 wire _2173_;
 wire _2174_;
 wire _2175_;
 wire _2176_;
 wire _2177_;
 wire _2178_;
 wire _2179_;
 wire _2180_;
 wire _2181_;
 wire _2182_;
 wire _2183_;
 wire _2184_;
 wire _2185_;
 wire _2186_;
 wire _2187_;
 wire _2188_;
 wire _2189_;
 wire _2190_;
 wire _2191_;
 wire _2192_;
 wire _2193_;
 wire _2194_;
 wire _2195_;
 wire _2196_;
 wire _2197_;
 wire _2198_;
 wire _2199_;
 wire _2200_;
 wire _2201_;
 wire _2202_;
 wire _2203_;
 wire _2204_;
 wire _2205_;
 wire _2206_;
 wire _2207_;
 wire _2208_;
 wire _2209_;
 wire _2210_;
 wire _2211_;
 wire _2212_;
 wire _2213_;
 wire _2214_;
 wire _2215_;
 wire _2216_;
 wire _2217_;
 wire _2218_;
 wire _2219_;
 wire _2220_;
 wire _2221_;
 wire _2222_;
 wire _2223_;
 wire _2224_;
 wire _2225_;
 wire _2226_;
 wire _2227_;
 wire _2228_;
 wire _2229_;
 wire _2230_;
 wire _2231_;
 wire _2232_;
 wire _2233_;
 wire _2234_;
 wire _2235_;
 wire _2236_;
 wire _2237_;
 wire _2238_;
 wire _2239_;
 wire _2240_;
 wire _2241_;
 wire _2242_;
 wire _2243_;
 wire _2244_;
 wire _2245_;
 wire _2246_;
 wire _2247_;
 wire _2248_;
 wire _2249_;
 wire _2250_;
 wire _2251_;
 wire _2252_;
 wire _2253_;
 wire _2254_;
 wire _2255_;
 wire _2256_;
 wire _2257_;
 wire _2258_;
 wire _2259_;
 wire _2260_;
 wire _2261_;
 wire _2262_;
 wire _2263_;
 wire _2264_;
 wire _2265_;
 wire _2266_;
 wire _2267_;
 wire _2268_;
 wire _2269_;
 wire _2270_;
 wire _2271_;
 wire _2272_;
 wire _2273_;
 wire _2274_;
 wire _2275_;
 wire _2276_;
 wire _2277_;
 wire _2278_;
 wire _2279_;
 wire _2280_;
 wire _2281_;
 wire _2282_;
 wire _2283_;
 wire _2284_;
 wire _2285_;
 wire _2286_;
 wire _2287_;
 wire _2288_;
 wire _2289_;
 wire _2290_;
 wire _2291_;
 wire _2292_;
 wire _2293_;
 wire _2294_;
 wire _2295_;
 wire _2296_;
 wire _2297_;
 wire _2298_;
 wire _2299_;
 wire _2300_;
 wire _2301_;
 wire _2302_;
 wire _2303_;
 wire _2304_;
 wire _2305_;
 wire _2306_;
 wire _2307_;
 wire _2308_;
 wire _2309_;
 wire _2310_;
 wire _2311_;
 wire _2312_;
 wire _2313_;
 wire _2314_;
 wire _2315_;
 wire _2316_;
 wire _2317_;
 wire _2318_;
 wire _2319_;
 wire _2320_;
 wire _2321_;
 wire _2322_;
 wire _2323_;
 wire _2324_;
 wire _2325_;
 wire _2326_;
 wire _2327_;
 wire _2328_;
 wire _2329_;
 wire _2330_;
 wire _2331_;
 wire _2332_;
 wire _2333_;
 wire _2334_;
 wire _2335_;
 wire _2336_;
 wire _2337_;
 wire _2338_;
 wire _2339_;
 wire _2340_;
 wire _2341_;
 wire _2342_;
 wire _2343_;
 wire _2344_;
 wire _2345_;
 wire _2346_;
 wire _2347_;
 wire _2348_;
 wire _2349_;
 wire _2350_;
 wire _2351_;
 wire _2352_;
 wire _2353_;
 wire _2354_;
 wire _2355_;
 wire _2356_;
 wire _2357_;
 wire _2358_;
 wire _2359_;
 wire _2360_;
 wire _2361_;
 wire _2362_;
 wire _2363_;
 wire _2364_;
 wire _2365_;
 wire _2366_;
 wire _2367_;
 wire _2368_;
 wire _2369_;
 wire _2370_;
 wire _2371_;
 wire _2372_;
 wire _2373_;
 wire _2374_;
 wire _2375_;
 wire _2376_;
 wire _2377_;
 wire _2378_;
 wire _2379_;
 wire _2380_;
 wire _2381_;
 wire _2382_;
 wire _2383_;
 wire _2384_;
 wire _2385_;
 wire _2386_;
 wire _2387_;
 wire _2388_;
 wire _2389_;
 wire _2390_;
 wire _2391_;
 wire _2392_;
 wire _2393_;
 wire _2394_;
 wire _2395_;
 wire _2396_;
 wire _2397_;
 wire _2398_;
 wire _2399_;
 wire _2400_;
 wire _2401_;
 wire _2402_;
 wire _2403_;
 wire _2404_;
 wire _2405_;
 wire _2406_;
 wire _2407_;
 wire _2408_;
 wire _2409_;
 wire _2410_;
 wire _2411_;
 wire _2412_;
 wire _2413_;
 wire _2414_;
 wire _2415_;
 wire _2416_;
 wire _2417_;
 wire _2418_;
 wire _2419_;
 wire _2420_;
 wire _2421_;
 wire _2422_;
 wire _2423_;
 wire _2424_;
 wire _2425_;
 wire _2426_;
 wire _2427_;
 wire _2428_;
 wire _2429_;
 wire _2430_;
 wire _2431_;
 wire _2432_;
 wire _2433_;
 wire _2434_;
 wire _2435_;
 wire _2436_;
 wire _2437_;
 wire _2438_;
 wire _2439_;
 wire _2440_;
 wire _2441_;
 wire _2442_;
 wire _2443_;
 wire _2444_;
 wire _2445_;
 wire _2446_;
 wire _2447_;
 wire _2448_;
 wire _2449_;
 wire _2450_;
 wire _2451_;
 wire _2452_;
 wire _2453_;
 wire _2454_;
 wire _2455_;
 wire _2456_;
 wire _2457_;
 wire _2458_;
 wire _2459_;
 wire _2460_;
 wire _2461_;
 wire _2462_;
 wire _2463_;
 wire _2464_;
 wire _2465_;
 wire _2466_;
 wire _2467_;
 wire _2468_;
 wire _2469_;
 wire _2470_;
 wire _2471_;
 wire _2472_;
 wire _2473_;
 wire _2474_;
 wire _2475_;
 wire _2476_;
 wire _2477_;
 wire _2478_;
 wire _2479_;
 wire _2480_;
 wire _2481_;
 wire _2482_;
 wire _2483_;
 wire _2484_;
 wire _2485_;
 wire _2486_;
 wire _2487_;
 wire _2488_;
 wire _2489_;
 wire _2490_;
 wire _2491_;
 wire _2492_;
 wire _2493_;
 wire _2494_;
 wire _2495_;
 wire _2496_;
 wire _2497_;
 wire _2498_;
 wire _2499_;
 wire _2500_;
 wire _2501_;
 wire _2502_;
 wire _2503_;
 wire _2504_;
 wire _2505_;
 wire _2506_;
 wire _2507_;
 wire _2508_;
 wire _2509_;
 wire _2510_;
 wire _2511_;
 wire _2512_;
 wire _2513_;
 wire _2514_;
 wire _2515_;
 wire _2516_;
 wire _2517_;
 wire _2518_;
 wire _2519_;
 wire _2520_;
 wire _2521_;
 wire _2522_;
 wire _2523_;
 wire _2524_;
 wire _2525_;
 wire _2526_;
 wire _2527_;
 wire _2528_;
 wire _2529_;
 wire _2530_;
 wire _2531_;
 wire _2532_;
 wire _2533_;
 wire _2534_;
 wire _2535_;
 wire _2536_;
 wire _2537_;
 wire _2538_;
 wire _2539_;
 wire _2540_;
 wire _2541_;
 wire _2542_;
 wire _2543_;
 wire _2544_;
 wire _2545_;
 wire _2546_;
 wire _2547_;
 wire _2548_;
 wire _2549_;
 wire _2550_;
 wire _2551_;
 wire _2552_;
 wire _2553_;
 wire _2554_;
 wire _2555_;
 wire _2556_;
 wire _2557_;
 wire _2558_;
 wire _2559_;
 wire _2560_;
 wire _2561_;
 wire _2562_;
 wire _2563_;
 wire _2564_;
 wire _2565_;
 wire _2566_;
 wire _2567_;
 wire _2568_;
 wire _2569_;
 wire _2570_;
 wire _2571_;
 wire _2572_;
 wire _2573_;
 wire _2574_;
 wire _2575_;
 wire _2576_;
 wire _2577_;
 wire _2578_;
 wire _2579_;
 wire _2580_;
 wire _2581_;
 wire _2582_;
 wire _2583_;
 wire _2584_;
 wire _2585_;
 wire _2586_;
 wire _2587_;
 wire _2588_;
 wire _2589_;
 wire _2590_;
 wire _2591_;
 wire _2592_;
 wire _2593_;
 wire _2594_;
 wire _2595_;
 wire _2596_;
 wire _2597_;
 wire _2598_;
 wire _2599_;
 wire _2600_;
 wire _2601_;
 wire _2602_;
 wire _2603_;
 wire _2604_;
 wire _2605_;
 wire _2606_;
 wire _2607_;
 wire _2608_;
 wire _2609_;
 wire _2610_;
 wire _2611_;
 wire _2612_;
 wire _2613_;
 wire _2614_;
 wire _2615_;
 wire _2616_;
 wire _2617_;
 wire _2618_;
 wire _2619_;
 wire _2620_;
 wire _2621_;
 wire _2622_;
 wire _2623_;
 wire _2624_;
 wire _2625_;
 wire _2626_;
 wire _2627_;
 wire _2628_;
 wire _2629_;
 wire _2630_;
 wire _2631_;
 wire _2632_;
 wire _2633_;
 wire _2634_;
 wire _2635_;
 wire _2636_;
 wire _2637_;
 wire _2638_;
 wire _2639_;
 wire _2640_;
 wire _2641_;
 wire _2642_;
 wire _2643_;
 wire _2644_;
 wire _2645_;
 wire _2646_;
 wire _2647_;
 wire _2648_;
 wire _2649_;
 wire _2650_;
 wire _2651_;
 wire _2652_;
 wire _2653_;
 wire _2654_;
 wire _2655_;
 wire _2656_;
 wire _2657_;
 wire _2658_;
 wire _2659_;
 wire _2660_;
 wire _2661_;
 wire _2662_;
 wire _2663_;
 wire _2664_;
 wire _2665_;
 wire _2666_;
 wire _2667_;
 wire _2668_;
 wire _2669_;
 wire _2670_;
 wire _2671_;
 wire _2672_;
 wire _2673_;
 wire _2674_;
 wire _2675_;
 wire _2676_;
 wire _2677_;
 wire _2678_;
 wire _2679_;
 wire _2680_;
 wire _2681_;
 wire _2682_;
 wire _2683_;
 wire _2684_;
 wire _2685_;
 wire _2686_;
 wire _2687_;
 wire _2688_;
 wire _2689_;
 wire _2690_;
 wire _2691_;
 wire _2692_;
 wire _2693_;
 wire _2694_;
 wire _2695_;
 wire _2696_;
 wire _2697_;
 wire _2698_;
 wire _2699_;
 wire _2700_;
 wire _2701_;
 wire _2702_;
 wire _2703_;
 wire _2704_;
 wire _2705_;
 wire _2706_;
 wire _2707_;
 wire _2708_;
 wire _2709_;
 wire _2710_;
 wire _2711_;
 wire _2712_;
 wire _2713_;
 wire _2714_;
 wire _2715_;
 wire _2716_;
 wire _2717_;
 wire _2718_;
 wire _2719_;
 wire _2720_;
 wire _2721_;
 wire _2722_;
 wire _2723_;
 wire _2724_;
 wire _2725_;
 wire _2726_;
 wire _2727_;
 wire _2728_;
 wire _2729_;
 wire _2730_;
 wire _2731_;
 wire _2732_;
 wire _2733_;
 wire _2734_;
 wire _2735_;
 wire _2736_;
 wire _2737_;
 wire _2738_;
 wire _2739_;
 wire _2740_;
 wire _2741_;
 wire _2742_;
 wire _2743_;
 wire _2744_;
 wire _2745_;
 wire _2746_;
 wire _2747_;
 wire _2748_;
 wire _2749_;
 wire _2750_;
 wire _2751_;
 wire _2752_;
 wire _2753_;
 wire _2754_;
 wire _2755_;
 wire _2756_;
 wire _2757_;
 wire _2758_;
 wire _2759_;
 wire _2760_;
 wire _2761_;
 wire _2762_;
 wire _2763_;
 wire _2764_;
 wire _2765_;
 wire _2766_;
 wire _2767_;
 wire _2768_;
 wire _2769_;
 wire _2770_;
 wire _2771_;
 wire _2772_;
 wire _2773_;
 wire _2774_;
 wire _2775_;
 wire _2776_;
 wire _2777_;
 wire _2778_;
 wire _2779_;
 wire _2780_;
 wire _2781_;
 wire _2782_;
 wire _2783_;
 wire _2784_;
 wire _2785_;
 wire _2786_;
 wire _2787_;
 wire _2788_;
 wire _2789_;
 wire _2790_;
 wire _2791_;
 wire _2792_;
 wire _2793_;
 wire _2794_;
 wire _2795_;
 wire _2796_;
 wire _2797_;
 wire _2798_;
 wire _2799_;
 wire _2800_;
 wire _2801_;
 wire _2802_;
 wire _2803_;
 wire _2804_;
 wire _2805_;
 wire _2806_;
 wire _2807_;
 wire _2808_;
 wire _2809_;
 wire _2810_;
 wire _2811_;
 wire _2812_;
 wire _2813_;
 wire _2814_;
 wire _2815_;
 wire _2816_;
 wire _2817_;
 wire _2818_;
 wire _2819_;
 wire _2820_;
 wire _2821_;
 wire _2822_;
 wire _2823_;
 wire _2824_;
 wire _2825_;
 wire _2826_;
 wire _2827_;
 wire _2828_;
 wire _2829_;
 wire _2830_;
 wire _2831_;
 wire _2832_;
 wire _2833_;
 wire _2834_;
 wire _2835_;
 wire _2836_;
 wire _2837_;
 wire _2838_;
 wire _2839_;
 wire _2840_;
 wire _2841_;
 wire _2842_;
 wire _2843_;
 wire _2844_;
 wire _2845_;
 wire _2846_;
 wire _2847_;
 wire _2848_;
 wire _2849_;
 wire _2850_;
 wire _2851_;
 wire _2852_;
 wire _2853_;
 wire _2854_;
 wire _2855_;
 wire _2856_;
 wire _2857_;
 wire _2858_;
 wire _2859_;
 wire _2860_;
 wire _2861_;
 wire _2862_;
 wire _2863_;
 wire _2864_;
 wire _2865_;
 wire _2866_;
 wire _2867_;
 wire _2868_;
 wire _2869_;
 wire _2870_;
 wire _2871_;
 wire _2872_;
 wire _2873_;
 wire _2874_;
 wire _2875_;
 wire _2876_;
 wire _2877_;
 wire _2878_;
 wire _2879_;
 wire _2880_;
 wire _2881_;
 wire _2882_;
 wire _2883_;
 wire _2884_;
 wire _2885_;
 wire _2886_;
 wire _2887_;
 wire _2888_;
 wire _2889_;
 wire _2890_;
 wire _2891_;
 wire _2892_;
 wire _2893_;
 wire _2894_;
 wire _2895_;
 wire _2896_;
 wire _2897_;
 wire _2898_;
 wire _2899_;
 wire _2900_;
 wire _2901_;
 wire _2902_;
 wire _2903_;
 wire _2904_;
 wire _2905_;
 wire _2906_;
 wire _2907_;
 wire _2908_;
 wire _2909_;
 wire _2910_;
 wire _2911_;
 wire _2912_;
 wire _2913_;
 wire _2914_;
 wire _2915_;
 wire _2916_;
 wire _2917_;
 wire _2918_;
 wire _2919_;
 wire _2920_;
 wire _2921_;
 wire _2922_;
 wire _2923_;
 wire _2924_;
 wire _2925_;
 wire _2926_;
 wire _2927_;
 wire _2928_;
 wire _2929_;
 wire _2930_;
 wire _2931_;
 wire _2932_;
 wire _2933_;
 wire _2934_;
 wire _2935_;
 wire _2936_;
 wire _2937_;
 wire _2938_;
 wire _2939_;
 wire _2940_;
 wire _2941_;
 wire _2942_;
 wire _2943_;
 wire _2944_;
 wire _2945_;
 wire _2946_;
 wire _2947_;
 wire _2948_;
 wire _2949_;
 wire _2950_;
 wire _2951_;
 wire _2952_;
 wire _2953_;
 wire _2954_;
 wire _2955_;
 wire _2956_;
 wire _2957_;
 wire _2958_;
 wire _2959_;
 wire _2960_;
 wire _2961_;
 wire _2962_;
 wire _2963_;
 wire _2964_;
 wire _2965_;
 wire _2966_;
 wire _2967_;
 wire _2968_;
 wire _2969_;
 wire _2970_;
 wire _2971_;
 wire _2972_;
 wire _2973_;
 wire _2974_;
 wire _2975_;
 wire _2976_;
 wire _2977_;
 wire _2978_;
 wire _2979_;
 wire _2980_;
 wire _2981_;
 wire _2982_;
 wire _2983_;
 wire _2984_;
 wire _2985_;
 wire _2986_;
 wire _2987_;
 wire _2988_;
 wire _2989_;
 wire _2990_;
 wire _2991_;
 wire _2992_;
 wire _2993_;
 wire _2994_;
 wire _2995_;
 wire _2996_;
 wire _2997_;
 wire _2998_;
 wire _2999_;
 wire _3000_;
 wire _3001_;
 wire _3002_;
 wire _3003_;
 wire _3004_;
 wire _3005_;
 wire _3006_;
 wire _3007_;
 wire _3008_;
 wire _3009_;
 wire _3010_;
 wire _3011_;
 wire _3012_;
 wire _3013_;
 wire _3014_;
 wire _3015_;
 wire _3016_;
 wire _3017_;
 wire _3018_;
 wire _3019_;
 wire _3020_;
 wire _3021_;
 wire _3022_;
 wire _3023_;
 wire _3024_;
 wire _3025_;
 wire _3026_;
 wire _3027_;
 wire _3028_;
 wire _3029_;
 wire _3030_;
 wire _3031_;
 wire _3032_;
 wire _3033_;
 wire _3034_;
 wire _3035_;
 wire _3036_;
 wire _3037_;
 wire _3038_;
 wire _3039_;
 wire _3040_;
 wire _3041_;
 wire _3042_;
 wire _3043_;
 wire _3044_;
 wire _3045_;
 wire _3046_;
 wire _3047_;
 wire _3048_;
 wire _3049_;
 wire _3050_;
 wire _3051_;
 wire _3052_;
 wire net93;
 wire net103;
 wire net104;
 wire net94;
 wire net105;
 wire net106;
 wire net226;
 wire net107;
 wire net108;
 wire net109;
 wire net95;
 wire net227;
 wire net228;
 wire net229;
 wire clknet_leaf_0_wb_clk_i;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net114;
 wire net115;
 wire net122;
 wire net116;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net131;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net132;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net133;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net134;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net135;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire \soc.boot_loading_offset[0] ;
 wire \soc.boot_loading_offset[1] ;
 wire \soc.boot_loading_offset[2] ;
 wire \soc.boot_loading_offset[3] ;
 wire \soc.boot_loading_offset[4] ;
 wire \soc.cpu.ALU.f ;
 wire \soc.cpu.ALU.no ;
 wire \soc.cpu.ALU.nx ;
 wire \soc.cpu.ALU.ny ;
 wire \soc.cpu.ALU.x[0] ;
 wire \soc.cpu.ALU.x[10] ;
 wire \soc.cpu.ALU.x[11] ;
 wire \soc.cpu.ALU.x[12] ;
 wire \soc.cpu.ALU.x[13] ;
 wire \soc.cpu.ALU.x[14] ;
 wire \soc.cpu.ALU.x[15] ;
 wire \soc.cpu.ALU.x[1] ;
 wire \soc.cpu.ALU.x[2] ;
 wire \soc.cpu.ALU.x[3] ;
 wire \soc.cpu.ALU.x[4] ;
 wire \soc.cpu.ALU.x[5] ;
 wire \soc.cpu.ALU.x[6] ;
 wire \soc.cpu.ALU.x[7] ;
 wire \soc.cpu.ALU.x[8] ;
 wire \soc.cpu.ALU.x[9] ;
 wire \soc.cpu.ALU.zx ;
 wire \soc.cpu.ALU.zy ;
 wire \soc.cpu.AReg.clk ;
 wire \soc.cpu.AReg.data[0] ;
 wire \soc.cpu.AReg.data[10] ;
 wire \soc.cpu.AReg.data[11] ;
 wire \soc.cpu.AReg.data[12] ;
 wire \soc.cpu.AReg.data[13] ;
 wire \soc.cpu.AReg.data[14] ;
 wire \soc.cpu.AReg.data[15] ;
 wire \soc.cpu.AReg.data[1] ;
 wire \soc.cpu.AReg.data[2] ;
 wire \soc.cpu.AReg.data[3] ;
 wire \soc.cpu.AReg.data[4] ;
 wire \soc.cpu.AReg.data[5] ;
 wire \soc.cpu.AReg.data[6] ;
 wire \soc.cpu.AReg.data[7] ;
 wire \soc.cpu.AReg.data[8] ;
 wire \soc.cpu.AReg.data[9] ;
 wire \soc.cpu.DMuxJMP.sel[0] ;
 wire \soc.cpu.DMuxJMP.sel[1] ;
 wire \soc.cpu.DMuxJMP.sel[2] ;
 wire \soc.cpu.PC.REG.data[0] ;
 wire \soc.cpu.PC.REG.data[10] ;
 wire \soc.cpu.PC.REG.data[11] ;
 wire \soc.cpu.PC.REG.data[12] ;
 wire \soc.cpu.PC.REG.data[13] ;
 wire \soc.cpu.PC.REG.data[14] ;
 wire \soc.cpu.PC.REG.data[1] ;
 wire \soc.cpu.PC.REG.data[2] ;
 wire \soc.cpu.PC.REG.data[3] ;
 wire \soc.cpu.PC.REG.data[4] ;
 wire \soc.cpu.PC.REG.data[5] ;
 wire \soc.cpu.PC.REG.data[6] ;
 wire \soc.cpu.PC.REG.data[7] ;
 wire \soc.cpu.PC.REG.data[8] ;
 wire \soc.cpu.PC.REG.data[9] ;
 wire \soc.cpu.PC.in[0] ;
 wire \soc.cpu.PC.in[10] ;
 wire \soc.cpu.PC.in[11] ;
 wire \soc.cpu.PC.in[12] ;
 wire \soc.cpu.PC.in[13] ;
 wire \soc.cpu.PC.in[14] ;
 wire \soc.cpu.PC.in[1] ;
 wire \soc.cpu.PC.in[2] ;
 wire \soc.cpu.PC.in[3] ;
 wire \soc.cpu.PC.in[4] ;
 wire \soc.cpu.PC.in[5] ;
 wire \soc.cpu.PC.in[6] ;
 wire \soc.cpu.PC.in[7] ;
 wire \soc.cpu.PC.in[8] ;
 wire \soc.cpu.PC.in[9] ;
 wire \soc.cpu.instruction[12] ;
 wire \soc.cpu.instruction[13] ;
 wire \soc.cpu.instruction[14] ;
 wire \soc.cpu.instruction[15] ;
 wire \soc.cpu.instruction[3] ;
 wire \soc.cpu.instruction[4] ;
 wire \soc.cpu.instruction[5] ;
 wire \soc.display_clks_before_active[0] ;
 wire \soc.gpio_i_stored[0] ;
 wire \soc.gpio_i_stored[1] ;
 wire \soc.gpio_i_stored[2] ;
 wire \soc.gpio_i_stored[3] ;
 wire \soc.hack_clk_strobe ;
 wire \soc.hack_clock_0.counter[0] ;
 wire \soc.hack_clock_0.counter[1] ;
 wire \soc.hack_clock_0.counter[2] ;
 wire \soc.hack_clock_0.counter[3] ;
 wire \soc.hack_clock_0.counter[4] ;
 wire \soc.hack_clock_0.counter[5] ;
 wire \soc.hack_clock_0.counter[6] ;
 wire \soc.hack_rom_request ;
 wire \soc.hack_wait_clocks[0] ;
 wire \soc.hack_wait_clocks[1] ;
 wire \soc.ram_data_out[0] ;
 wire \soc.ram_data_out[10] ;
 wire \soc.ram_data_out[11] ;
 wire \soc.ram_data_out[12] ;
 wire \soc.ram_data_out[13] ;
 wire \soc.ram_data_out[14] ;
 wire \soc.ram_data_out[15] ;
 wire \soc.ram_data_out[1] ;
 wire \soc.ram_data_out[2] ;
 wire \soc.ram_data_out[3] ;
 wire \soc.ram_data_out[4] ;
 wire \soc.ram_data_out[5] ;
 wire \soc.ram_data_out[6] ;
 wire \soc.ram_data_out[7] ;
 wire \soc.ram_data_out[8] ;
 wire \soc.ram_data_out[9] ;
 wire \soc.ram_encoder_0.address[0] ;
 wire \soc.ram_encoder_0.address[10] ;
 wire \soc.ram_encoder_0.address[11] ;
 wire \soc.ram_encoder_0.address[12] ;
 wire \soc.ram_encoder_0.address[13] ;
 wire \soc.ram_encoder_0.address[14] ;
 wire \soc.ram_encoder_0.address[1] ;
 wire \soc.ram_encoder_0.address[2] ;
 wire \soc.ram_encoder_0.address[3] ;
 wire \soc.ram_encoder_0.address[4] ;
 wire \soc.ram_encoder_0.address[5] ;
 wire \soc.ram_encoder_0.address[6] ;
 wire \soc.ram_encoder_0.address[7] ;
 wire \soc.ram_encoder_0.address[8] ;
 wire \soc.ram_encoder_0.address[9] ;
 wire \soc.ram_encoder_0.current_state[0] ;
 wire \soc.ram_encoder_0.current_state[1] ;
 wire \soc.ram_encoder_0.current_state[2] ;
 wire \soc.ram_encoder_0.data_out[0] ;
 wire \soc.ram_encoder_0.data_out[10] ;
 wire \soc.ram_encoder_0.data_out[11] ;
 wire \soc.ram_encoder_0.data_out[12] ;
 wire \soc.ram_encoder_0.data_out[13] ;
 wire \soc.ram_encoder_0.data_out[14] ;
 wire \soc.ram_encoder_0.data_out[15] ;
 wire \soc.ram_encoder_0.data_out[1] ;
 wire \soc.ram_encoder_0.data_out[2] ;
 wire \soc.ram_encoder_0.data_out[3] ;
 wire \soc.ram_encoder_0.data_out[4] ;
 wire \soc.ram_encoder_0.data_out[5] ;
 wire \soc.ram_encoder_0.data_out[6] ;
 wire \soc.ram_encoder_0.data_out[7] ;
 wire \soc.ram_encoder_0.data_out[8] ;
 wire \soc.ram_encoder_0.data_out[9] ;
 wire \soc.ram_encoder_0.initialized ;
 wire \soc.ram_encoder_0.initializing_step[0] ;
 wire \soc.ram_encoder_0.initializing_step[1] ;
 wire \soc.ram_encoder_0.initializing_step[2] ;
 wire \soc.ram_encoder_0.initializing_step[3] ;
 wire \soc.ram_encoder_0.initializing_step[4] ;
 wire \soc.ram_encoder_0.input_bits_left[2] ;
 wire \soc.ram_encoder_0.input_bits_left[3] ;
 wire \soc.ram_encoder_0.input_bits_left[4] ;
 wire \soc.ram_encoder_0.input_buffer[0] ;
 wire \soc.ram_encoder_0.input_buffer[10] ;
 wire \soc.ram_encoder_0.input_buffer[11] ;
 wire \soc.ram_encoder_0.input_buffer[1] ;
 wire \soc.ram_encoder_0.input_buffer[2] ;
 wire \soc.ram_encoder_0.input_buffer[3] ;
 wire \soc.ram_encoder_0.input_buffer[4] ;
 wire \soc.ram_encoder_0.input_buffer[5] ;
 wire \soc.ram_encoder_0.input_buffer[6] ;
 wire \soc.ram_encoder_0.input_buffer[7] ;
 wire \soc.ram_encoder_0.input_buffer[8] ;
 wire \soc.ram_encoder_0.input_buffer[9] ;
 wire \soc.ram_encoder_0.output_bits_left[2] ;
 wire \soc.ram_encoder_0.output_bits_left[3] ;
 wire \soc.ram_encoder_0.output_bits_left[4] ;
 wire \soc.ram_encoder_0.output_buffer[10] ;
 wire \soc.ram_encoder_0.output_buffer[11] ;
 wire \soc.ram_encoder_0.output_buffer[12] ;
 wire \soc.ram_encoder_0.output_buffer[13] ;
 wire \soc.ram_encoder_0.output_buffer[14] ;
 wire \soc.ram_encoder_0.output_buffer[15] ;
 wire \soc.ram_encoder_0.output_buffer[16] ;
 wire \soc.ram_encoder_0.output_buffer[17] ;
 wire \soc.ram_encoder_0.output_buffer[18] ;
 wire \soc.ram_encoder_0.output_buffer[19] ;
 wire \soc.ram_encoder_0.output_buffer[1] ;
 wire \soc.ram_encoder_0.output_buffer[2] ;
 wire \soc.ram_encoder_0.output_buffer[3] ;
 wire \soc.ram_encoder_0.output_buffer[4] ;
 wire \soc.ram_encoder_0.output_buffer[5] ;
 wire \soc.ram_encoder_0.output_buffer[6] ;
 wire \soc.ram_encoder_0.output_buffer[7] ;
 wire \soc.ram_encoder_0.output_buffer[8] ;
 wire \soc.ram_encoder_0.output_buffer[9] ;
 wire \soc.ram_encoder_0.request_address[0] ;
 wire \soc.ram_encoder_0.request_address[10] ;
 wire \soc.ram_encoder_0.request_address[11] ;
 wire \soc.ram_encoder_0.request_address[12] ;
 wire \soc.ram_encoder_0.request_address[13] ;
 wire \soc.ram_encoder_0.request_address[14] ;
 wire \soc.ram_encoder_0.request_address[1] ;
 wire \soc.ram_encoder_0.request_address[2] ;
 wire \soc.ram_encoder_0.request_address[3] ;
 wire \soc.ram_encoder_0.request_address[4] ;
 wire \soc.ram_encoder_0.request_address[5] ;
 wire \soc.ram_encoder_0.request_address[6] ;
 wire \soc.ram_encoder_0.request_address[7] ;
 wire \soc.ram_encoder_0.request_address[8] ;
 wire \soc.ram_encoder_0.request_address[9] ;
 wire \soc.ram_encoder_0.request_data_out[0] ;
 wire \soc.ram_encoder_0.request_data_out[10] ;
 wire \soc.ram_encoder_0.request_data_out[11] ;
 wire \soc.ram_encoder_0.request_data_out[12] ;
 wire \soc.ram_encoder_0.request_data_out[13] ;
 wire \soc.ram_encoder_0.request_data_out[14] ;
 wire \soc.ram_encoder_0.request_data_out[15] ;
 wire \soc.ram_encoder_0.request_data_out[1] ;
 wire \soc.ram_encoder_0.request_data_out[2] ;
 wire \soc.ram_encoder_0.request_data_out[3] ;
 wire \soc.ram_encoder_0.request_data_out[4] ;
 wire \soc.ram_encoder_0.request_data_out[5] ;
 wire \soc.ram_encoder_0.request_data_out[6] ;
 wire \soc.ram_encoder_0.request_data_out[7] ;
 wire \soc.ram_encoder_0.request_data_out[8] ;
 wire \soc.ram_encoder_0.request_data_out[9] ;
 wire \soc.ram_encoder_0.request_write ;
 wire \soc.ram_encoder_0.sram_sio_oe ;
 wire \soc.ram_encoder_0.toggled_sram_sck ;
 wire \soc.ram_step1_write_request ;
 wire \soc.ram_step2_read_request ;
 wire \soc.rom_encoder_0.current_state[0] ;
 wire \soc.rom_encoder_0.current_state[1] ;
 wire \soc.rom_encoder_0.current_state[2] ;
 wire \soc.rom_encoder_0.data_out[0] ;
 wire \soc.rom_encoder_0.data_out[10] ;
 wire \soc.rom_encoder_0.data_out[11] ;
 wire \soc.rom_encoder_0.data_out[12] ;
 wire \soc.rom_encoder_0.data_out[13] ;
 wire \soc.rom_encoder_0.data_out[14] ;
 wire \soc.rom_encoder_0.data_out[15] ;
 wire \soc.rom_encoder_0.data_out[1] ;
 wire \soc.rom_encoder_0.data_out[2] ;
 wire \soc.rom_encoder_0.data_out[3] ;
 wire \soc.rom_encoder_0.data_out[4] ;
 wire \soc.rom_encoder_0.data_out[5] ;
 wire \soc.rom_encoder_0.data_out[6] ;
 wire \soc.rom_encoder_0.data_out[7] ;
 wire \soc.rom_encoder_0.data_out[8] ;
 wire \soc.rom_encoder_0.data_out[9] ;
 wire \soc.rom_encoder_0.initialized ;
 wire \soc.rom_encoder_0.initializing_step[0] ;
 wire \soc.rom_encoder_0.initializing_step[1] ;
 wire \soc.rom_encoder_0.initializing_step[2] ;
 wire \soc.rom_encoder_0.initializing_step[3] ;
 wire \soc.rom_encoder_0.initializing_step[4] ;
 wire \soc.rom_encoder_0.input_bits_left[2] ;
 wire \soc.rom_encoder_0.input_bits_left[3] ;
 wire \soc.rom_encoder_0.input_bits_left[4] ;
 wire \soc.rom_encoder_0.input_buffer[0] ;
 wire \soc.rom_encoder_0.input_buffer[10] ;
 wire \soc.rom_encoder_0.input_buffer[11] ;
 wire \soc.rom_encoder_0.input_buffer[1] ;
 wire \soc.rom_encoder_0.input_buffer[2] ;
 wire \soc.rom_encoder_0.input_buffer[3] ;
 wire \soc.rom_encoder_0.input_buffer[4] ;
 wire \soc.rom_encoder_0.input_buffer[5] ;
 wire \soc.rom_encoder_0.input_buffer[6] ;
 wire \soc.rom_encoder_0.input_buffer[7] ;
 wire \soc.rom_encoder_0.input_buffer[8] ;
 wire \soc.rom_encoder_0.input_buffer[9] ;
 wire \soc.rom_encoder_0.output_bits_left[2] ;
 wire \soc.rom_encoder_0.output_bits_left[3] ;
 wire \soc.rom_encoder_0.output_bits_left[4] ;
 wire \soc.rom_encoder_0.output_buffer[10] ;
 wire \soc.rom_encoder_0.output_buffer[11] ;
 wire \soc.rom_encoder_0.output_buffer[12] ;
 wire \soc.rom_encoder_0.output_buffer[13] ;
 wire \soc.rom_encoder_0.output_buffer[14] ;
 wire \soc.rom_encoder_0.output_buffer[15] ;
 wire \soc.rom_encoder_0.output_buffer[16] ;
 wire \soc.rom_encoder_0.output_buffer[17] ;
 wire \soc.rom_encoder_0.output_buffer[18] ;
 wire \soc.rom_encoder_0.output_buffer[19] ;
 wire \soc.rom_encoder_0.output_buffer[1] ;
 wire \soc.rom_encoder_0.output_buffer[2] ;
 wire \soc.rom_encoder_0.output_buffer[3] ;
 wire \soc.rom_encoder_0.output_buffer[4] ;
 wire \soc.rom_encoder_0.output_buffer[5] ;
 wire \soc.rom_encoder_0.output_buffer[6] ;
 wire \soc.rom_encoder_0.output_buffer[7] ;
 wire \soc.rom_encoder_0.output_buffer[8] ;
 wire \soc.rom_encoder_0.output_buffer[9] ;
 wire \soc.rom_encoder_0.request_address[0] ;
 wire \soc.rom_encoder_0.request_address[10] ;
 wire \soc.rom_encoder_0.request_address[11] ;
 wire \soc.rom_encoder_0.request_address[12] ;
 wire \soc.rom_encoder_0.request_address[13] ;
 wire \soc.rom_encoder_0.request_address[14] ;
 wire \soc.rom_encoder_0.request_address[1] ;
 wire \soc.rom_encoder_0.request_address[2] ;
 wire \soc.rom_encoder_0.request_address[3] ;
 wire \soc.rom_encoder_0.request_address[4] ;
 wire \soc.rom_encoder_0.request_address[5] ;
 wire \soc.rom_encoder_0.request_address[6] ;
 wire \soc.rom_encoder_0.request_address[7] ;
 wire \soc.rom_encoder_0.request_address[8] ;
 wire \soc.rom_encoder_0.request_address[9] ;
 wire \soc.rom_encoder_0.request_data_out[0] ;
 wire \soc.rom_encoder_0.request_data_out[10] ;
 wire \soc.rom_encoder_0.request_data_out[11] ;
 wire \soc.rom_encoder_0.request_data_out[12] ;
 wire \soc.rom_encoder_0.request_data_out[13] ;
 wire \soc.rom_encoder_0.request_data_out[14] ;
 wire \soc.rom_encoder_0.request_data_out[15] ;
 wire \soc.rom_encoder_0.request_data_out[1] ;
 wire \soc.rom_encoder_0.request_data_out[2] ;
 wire \soc.rom_encoder_0.request_data_out[3] ;
 wire \soc.rom_encoder_0.request_data_out[4] ;
 wire \soc.rom_encoder_0.request_data_out[5] ;
 wire \soc.rom_encoder_0.request_data_out[6] ;
 wire \soc.rom_encoder_0.request_data_out[7] ;
 wire \soc.rom_encoder_0.request_data_out[8] ;
 wire \soc.rom_encoder_0.request_data_out[9] ;
 wire \soc.rom_encoder_0.request_write ;
 wire \soc.rom_encoder_0.sram_sio_oe ;
 wire \soc.rom_encoder_0.toggled_sram_sck ;
 wire \soc.rom_encoder_0.write_enable ;
 wire \soc.rom_loader.current_address[0] ;
 wire \soc.rom_loader.current_address[10] ;
 wire \soc.rom_loader.current_address[11] ;
 wire \soc.rom_loader.current_address[12] ;
 wire \soc.rom_loader.current_address[13] ;
 wire \soc.rom_loader.current_address[14] ;
 wire \soc.rom_loader.current_address[1] ;
 wire \soc.rom_loader.current_address[2] ;
 wire \soc.rom_loader.current_address[3] ;
 wire \soc.rom_loader.current_address[4] ;
 wire \soc.rom_loader.current_address[5] ;
 wire \soc.rom_loader.current_address[6] ;
 wire \soc.rom_loader.current_address[7] ;
 wire \soc.rom_loader.current_address[8] ;
 wire \soc.rom_loader.current_address[9] ;
 wire \soc.rom_loader.rom_request ;
 wire \soc.rom_loader.wait_fall_clk ;
 wire \soc.rom_loader.was_loading ;
 wire \soc.rom_loader.writing ;
 wire \soc.spi_video_ram_1.buffer_index[0] ;
 wire \soc.spi_video_ram_1.buffer_index[1] ;
 wire \soc.spi_video_ram_1.buffer_index[2] ;
 wire \soc.spi_video_ram_1.buffer_index[3] ;
 wire \soc.spi_video_ram_1.buffer_index[4] ;
 wire \soc.spi_video_ram_1.buffer_index[5] ;
 wire \soc.spi_video_ram_1.current_state[0] ;
 wire \soc.spi_video_ram_1.current_state[1] ;
 wire \soc.spi_video_ram_1.current_state[2] ;
 wire \soc.spi_video_ram_1.current_state[3] ;
 wire \soc.spi_video_ram_1.current_state[4] ;
 wire \soc.spi_video_ram_1.fifo_in_address[0] ;
 wire \soc.spi_video_ram_1.fifo_in_address[10] ;
 wire \soc.spi_video_ram_1.fifo_in_address[11] ;
 wire \soc.spi_video_ram_1.fifo_in_address[12] ;
 wire \soc.spi_video_ram_1.fifo_in_address[1] ;
 wire \soc.spi_video_ram_1.fifo_in_address[2] ;
 wire \soc.spi_video_ram_1.fifo_in_address[3] ;
 wire \soc.spi_video_ram_1.fifo_in_address[4] ;
 wire \soc.spi_video_ram_1.fifo_in_address[5] ;
 wire \soc.spi_video_ram_1.fifo_in_address[6] ;
 wire \soc.spi_video_ram_1.fifo_in_address[7] ;
 wire \soc.spi_video_ram_1.fifo_in_address[8] ;
 wire \soc.spi_video_ram_1.fifo_in_address[9] ;
 wire \soc.spi_video_ram_1.fifo_in_data[0] ;
 wire \soc.spi_video_ram_1.fifo_in_data[10] ;
 wire \soc.spi_video_ram_1.fifo_in_data[11] ;
 wire \soc.spi_video_ram_1.fifo_in_data[12] ;
 wire \soc.spi_video_ram_1.fifo_in_data[13] ;
 wire \soc.spi_video_ram_1.fifo_in_data[14] ;
 wire \soc.spi_video_ram_1.fifo_in_data[15] ;
 wire \soc.spi_video_ram_1.fifo_in_data[1] ;
 wire \soc.spi_video_ram_1.fifo_in_data[2] ;
 wire \soc.spi_video_ram_1.fifo_in_data[3] ;
 wire \soc.spi_video_ram_1.fifo_in_data[4] ;
 wire \soc.spi_video_ram_1.fifo_in_data[5] ;
 wire \soc.spi_video_ram_1.fifo_in_data[6] ;
 wire \soc.spi_video_ram_1.fifo_in_data[7] ;
 wire \soc.spi_video_ram_1.fifo_in_data[8] ;
 wire \soc.spi_video_ram_1.fifo_in_data[9] ;
 wire \soc.spi_video_ram_1.fifo_read_request ;
 wire \soc.spi_video_ram_1.fifo_write_request ;
 wire \soc.spi_video_ram_1.initialized ;
 wire \soc.spi_video_ram_1.output_buffer[10] ;
 wire \soc.spi_video_ram_1.output_buffer[11] ;
 wire \soc.spi_video_ram_1.output_buffer[12] ;
 wire \soc.spi_video_ram_1.output_buffer[13] ;
 wire \soc.spi_video_ram_1.output_buffer[14] ;
 wire \soc.spi_video_ram_1.output_buffer[15] ;
 wire \soc.spi_video_ram_1.output_buffer[16] ;
 wire \soc.spi_video_ram_1.output_buffer[17] ;
 wire \soc.spi_video_ram_1.output_buffer[18] ;
 wire \soc.spi_video_ram_1.output_buffer[19] ;
 wire \soc.spi_video_ram_1.output_buffer[1] ;
 wire \soc.spi_video_ram_1.output_buffer[20] ;
 wire \soc.spi_video_ram_1.output_buffer[21] ;
 wire \soc.spi_video_ram_1.output_buffer[22] ;
 wire \soc.spi_video_ram_1.output_buffer[23] ;
 wire \soc.spi_video_ram_1.output_buffer[2] ;
 wire \soc.spi_video_ram_1.output_buffer[3] ;
 wire \soc.spi_video_ram_1.output_buffer[4] ;
 wire \soc.spi_video_ram_1.output_buffer[5] ;
 wire \soc.spi_video_ram_1.output_buffer[6] ;
 wire \soc.spi_video_ram_1.output_buffer[7] ;
 wire \soc.spi_video_ram_1.output_buffer[8] ;
 wire \soc.spi_video_ram_1.output_buffer[9] ;
 wire \soc.spi_video_ram_1.read_value[0] ;
 wire \soc.spi_video_ram_1.read_value[1] ;
 wire \soc.spi_video_ram_1.read_value[2] ;
 wire \soc.spi_video_ram_1.read_value[3] ;
 wire \soc.spi_video_ram_1.sram_sck_fall_edge ;
 wire \soc.spi_video_ram_1.sram_sck_rise_edge ;
 wire \soc.spi_video_ram_1.sram_sio_oe ;
 wire \soc.spi_video_ram_1.start_read ;
 wire \soc.spi_video_ram_1.state_counter[0] ;
 wire \soc.spi_video_ram_1.state_counter[10] ;
 wire \soc.spi_video_ram_1.state_counter[1] ;
 wire \soc.spi_video_ram_1.state_counter[2] ;
 wire \soc.spi_video_ram_1.state_counter[3] ;
 wire \soc.spi_video_ram_1.state_counter[4] ;
 wire \soc.spi_video_ram_1.state_counter[5] ;
 wire \soc.spi_video_ram_1.state_counter[6] ;
 wire \soc.spi_video_ram_1.state_counter[7] ;
 wire \soc.spi_video_ram_1.state_counter[8] ;
 wire \soc.spi_video_ram_1.state_counter[9] ;
 wire \soc.spi_video_ram_1.state_sram_clk_counter[0] ;
 wire \soc.spi_video_ram_1.state_sram_clk_counter[1] ;
 wire \soc.spi_video_ram_1.state_sram_clk_counter[2] ;
 wire \soc.spi_video_ram_1.state_sram_clk_counter[3] ;
 wire \soc.spi_video_ram_1.state_sram_clk_counter[4] ;
 wire \soc.spi_video_ram_1.state_sram_clk_counter[5] ;
 wire \soc.spi_video_ram_1.state_sram_clk_counter[6] ;
 wire \soc.spi_video_ram_1.state_sram_clk_counter[7] ;
 wire \soc.spi_video_ram_1.state_sram_clk_counter[8] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[0][0] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[0][10] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[0][11] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[0][12] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[0][13] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[0][14] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[0][15] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[0][16] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[0][17] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[0][18] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[0][19] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[0][1] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[0][20] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[0][21] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[0][22] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[0][23] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[0][24] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[0][25] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[0][26] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[0][27] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[0][28] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[0][2] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[0][3] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[0][4] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[0][5] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[0][6] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[0][7] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[0][8] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[0][9] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[1][0] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[1][10] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[1][11] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[1][12] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[1][13] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[1][14] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[1][15] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[1][16] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[1][17] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[1][18] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[1][19] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[1][1] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[1][20] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[1][21] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[1][22] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[1][23] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[1][24] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[1][25] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[1][26] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[1][27] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[1][28] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[1][2] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[1][3] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[1][4] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[1][5] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[1][6] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[1][7] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[1][8] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[1][9] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[2][0] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[2][10] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[2][11] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[2][12] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[2][13] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[2][14] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[2][15] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[2][16] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[2][17] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[2][18] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[2][19] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[2][1] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[2][20] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[2][21] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[2][22] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[2][23] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[2][24] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[2][25] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[2][26] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[2][27] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[2][28] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[2][2] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[2][3] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[2][4] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[2][5] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[2][6] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[2][7] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[2][8] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[2][9] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[3][0] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[3][10] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[3][11] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[3][12] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[3][13] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[3][14] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[3][15] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[3][16] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[3][17] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[3][18] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[3][19] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[3][1] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[3][20] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[3][21] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[3][22] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[3][23] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[3][24] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[3][25] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[3][26] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[3][27] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[3][28] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[3][2] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[3][3] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[3][4] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[3][5] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[3][6] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[3][7] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[3][8] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[3][9] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[4][0] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[4][10] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[4][11] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[4][12] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[4][13] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[4][14] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[4][15] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[4][16] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[4][17] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[4][18] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[4][19] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[4][1] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[4][20] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[4][21] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[4][22] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[4][23] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[4][24] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[4][25] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[4][26] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[4][27] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[4][28] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[4][2] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[4][3] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[4][4] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[4][5] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[4][6] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[4][7] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[4][8] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[4][9] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[5][0] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[5][10] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[5][11] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[5][12] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[5][13] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[5][14] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[5][15] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[5][16] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[5][17] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[5][18] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[5][19] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[5][1] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[5][20] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[5][21] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[5][22] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[5][23] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[5][24] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[5][25] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[5][26] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[5][27] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[5][28] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[5][2] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[5][3] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[5][4] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[5][5] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[5][6] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[5][7] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[5][8] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[5][9] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[6][0] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[6][10] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[6][11] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[6][12] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[6][13] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[6][14] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[6][15] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[6][16] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[6][17] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[6][18] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[6][19] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[6][1] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[6][20] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[6][21] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[6][22] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[6][23] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[6][24] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[6][25] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[6][26] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[6][27] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[6][28] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[6][2] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[6][3] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[6][4] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[6][5] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[6][6] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[6][7] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[6][8] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[6][9] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[7][0] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[7][10] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[7][11] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[7][12] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[7][13] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[7][14] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[7][15] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[7][16] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[7][17] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[7][18] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[7][19] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[7][1] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[7][20] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[7][21] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[7][22] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[7][23] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[7][24] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[7][25] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[7][26] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[7][27] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[7][28] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[7][2] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[7][3] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[7][4] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[7][5] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[7][6] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[7][7] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[7][8] ;
 wire \soc.spi_video_ram_1.write_fifo.fifo_mem[7][9] ;
 wire \soc.spi_video_ram_1.write_fifo.read_pointer[0] ;
 wire \soc.spi_video_ram_1.write_fifo.read_pointer[1] ;
 wire \soc.spi_video_ram_1.write_fifo.read_pointer[2] ;
 wire \soc.spi_video_ram_1.write_fifo.write_pointer[0] ;
 wire \soc.spi_video_ram_1.write_fifo.write_pointer[1] ;
 wire \soc.spi_video_ram_1.write_fifo.write_pointer[2] ;
 wire \soc.synch_hack_writeM ;
 wire \soc.video_generator_1.h_count[1] ;
 wire \soc.video_generator_1.h_count[2] ;
 wire \soc.video_generator_1.h_count[3] ;
 wire \soc.video_generator_1.h_count[4] ;
 wire \soc.video_generator_1.h_count[5] ;
 wire \soc.video_generator_1.h_count[6] ;
 wire \soc.video_generator_1.h_count[7] ;
 wire \soc.video_generator_1.h_count[8] ;
 wire \soc.video_generator_1.h_count[9] ;
 wire \soc.video_generator_1.v_count[0] ;
 wire \soc.video_generator_1.v_count[1] ;
 wire \soc.video_generator_1.v_count[2] ;
 wire \soc.video_generator_1.v_count[3] ;
 wire \soc.video_generator_1.v_count[4] ;
 wire \soc.video_generator_1.v_count[5] ;
 wire \soc.video_generator_1.v_count[6] ;
 wire \soc.video_generator_1.v_count[7] ;
 wire \soc.video_generator_1.v_count[8] ;
 wire \soc.video_generator_1.v_count[9] ;
 wire net193;
 wire net194;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net195;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net196;
 wire net224;
 wire net225;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire clknet_leaf_1_wb_clk_i;
 wire clknet_leaf_2_wb_clk_i;
 wire clknet_leaf_3_wb_clk_i;
 wire clknet_leaf_4_wb_clk_i;
 wire clknet_leaf_5_wb_clk_i;
 wire clknet_leaf_6_wb_clk_i;
 wire clknet_leaf_7_wb_clk_i;
 wire clknet_leaf_8_wb_clk_i;
 wire clknet_leaf_9_wb_clk_i;
 wire clknet_leaf_10_wb_clk_i;
 wire clknet_leaf_11_wb_clk_i;
 wire clknet_leaf_12_wb_clk_i;
 wire clknet_leaf_13_wb_clk_i;
 wire clknet_leaf_14_wb_clk_i;
 wire clknet_leaf_15_wb_clk_i;
 wire clknet_leaf_16_wb_clk_i;
 wire clknet_leaf_17_wb_clk_i;
 wire clknet_leaf_18_wb_clk_i;
 wire clknet_leaf_19_wb_clk_i;
 wire clknet_leaf_20_wb_clk_i;
 wire clknet_leaf_21_wb_clk_i;
 wire clknet_leaf_22_wb_clk_i;
 wire clknet_leaf_23_wb_clk_i;
 wire clknet_leaf_24_wb_clk_i;
 wire clknet_leaf_25_wb_clk_i;
 wire clknet_leaf_26_wb_clk_i;
 wire clknet_leaf_27_wb_clk_i;
 wire clknet_leaf_28_wb_clk_i;
 wire clknet_leaf_29_wb_clk_i;
 wire clknet_leaf_30_wb_clk_i;
 wire clknet_leaf_31_wb_clk_i;
 wire clknet_leaf_32_wb_clk_i;
 wire clknet_leaf_33_wb_clk_i;
 wire clknet_leaf_34_wb_clk_i;
 wire clknet_leaf_35_wb_clk_i;
 wire clknet_leaf_36_wb_clk_i;
 wire clknet_leaf_37_wb_clk_i;
 wire clknet_leaf_38_wb_clk_i;
 wire clknet_leaf_39_wb_clk_i;
 wire clknet_leaf_40_wb_clk_i;
 wire clknet_leaf_41_wb_clk_i;
 wire clknet_leaf_42_wb_clk_i;
 wire clknet_leaf_43_wb_clk_i;
 wire clknet_leaf_44_wb_clk_i;
 wire clknet_leaf_45_wb_clk_i;
 wire clknet_leaf_46_wb_clk_i;
 wire clknet_leaf_47_wb_clk_i;
 wire clknet_leaf_48_wb_clk_i;
 wire clknet_leaf_49_wb_clk_i;
 wire clknet_leaf_50_wb_clk_i;
 wire clknet_leaf_51_wb_clk_i;
 wire clknet_leaf_52_wb_clk_i;
 wire clknet_leaf_53_wb_clk_i;
 wire clknet_leaf_54_wb_clk_i;
 wire clknet_leaf_55_wb_clk_i;
 wire clknet_leaf_56_wb_clk_i;
 wire clknet_leaf_57_wb_clk_i;
 wire clknet_leaf_58_wb_clk_i;
 wire clknet_leaf_59_wb_clk_i;
 wire clknet_leaf_60_wb_clk_i;
 wire clknet_leaf_61_wb_clk_i;
 wire clknet_leaf_62_wb_clk_i;
 wire clknet_leaf_63_wb_clk_i;
 wire clknet_leaf_64_wb_clk_i;
 wire clknet_leaf_65_wb_clk_i;
 wire clknet_leaf_66_wb_clk_i;
 wire clknet_leaf_67_wb_clk_i;
 wire clknet_leaf_70_wb_clk_i;
 wire clknet_leaf_72_wb_clk_i;
 wire clknet_leaf_73_wb_clk_i;
 wire clknet_leaf_74_wb_clk_i;
 wire clknet_leaf_75_wb_clk_i;
 wire clknet_leaf_76_wb_clk_i;
 wire clknet_leaf_77_wb_clk_i;
 wire clknet_leaf_78_wb_clk_i;
 wire clknet_leaf_79_wb_clk_i;
 wire clknet_leaf_80_wb_clk_i;
 wire clknet_leaf_81_wb_clk_i;
 wire clknet_leaf_82_wb_clk_i;
 wire clknet_leaf_83_wb_clk_i;
 wire clknet_leaf_84_wb_clk_i;
 wire clknet_leaf_85_wb_clk_i;
 wire clknet_leaf_86_wb_clk_i;
 wire clknet_leaf_87_wb_clk_i;
 wire clknet_leaf_88_wb_clk_i;
 wire clknet_leaf_89_wb_clk_i;
 wire clknet_leaf_90_wb_clk_i;
 wire clknet_leaf_91_wb_clk_i;
 wire clknet_leaf_92_wb_clk_i;
 wire clknet_leaf_93_wb_clk_i;
 wire clknet_leaf_94_wb_clk_i;
 wire clknet_leaf_95_wb_clk_i;
 wire clknet_leaf_96_wb_clk_i;
 wire clknet_leaf_97_wb_clk_i;
 wire clknet_leaf_98_wb_clk_i;
 wire clknet_leaf_99_wb_clk_i;
 wire clknet_leaf_100_wb_clk_i;
 wire clknet_leaf_101_wb_clk_i;
 wire clknet_leaf_103_wb_clk_i;
 wire clknet_leaf_104_wb_clk_i;
 wire clknet_leaf_105_wb_clk_i;
 wire clknet_leaf_106_wb_clk_i;
 wire clknet_leaf_107_wb_clk_i;
 wire clknet_leaf_108_wb_clk_i;
 wire clknet_leaf_109_wb_clk_i;
 wire clknet_leaf_110_wb_clk_i;
 wire clknet_leaf_111_wb_clk_i;
 wire clknet_leaf_112_wb_clk_i;
 wire clknet_leaf_113_wb_clk_i;
 wire clknet_leaf_114_wb_clk_i;
 wire clknet_leaf_115_wb_clk_i;
 wire clknet_leaf_116_wb_clk_i;
 wire clknet_leaf_117_wb_clk_i;
 wire clknet_leaf_118_wb_clk_i;
 wire clknet_leaf_119_wb_clk_i;
 wire clknet_leaf_120_wb_clk_i;
 wire clknet_leaf_121_wb_clk_i;
 wire clknet_leaf_122_wb_clk_i;
 wire clknet_leaf_123_wb_clk_i;
 wire clknet_leaf_124_wb_clk_i;
 wire clknet_leaf_125_wb_clk_i;
 wire clknet_leaf_126_wb_clk_i;
 wire clknet_leaf_127_wb_clk_i;
 wire clknet_leaf_128_wb_clk_i;
 wire clknet_leaf_129_wb_clk_i;
 wire clknet_leaf_130_wb_clk_i;
 wire clknet_leaf_131_wb_clk_i;
 wire clknet_leaf_132_wb_clk_i;
 wire clknet_leaf_133_wb_clk_i;
 wire clknet_leaf_134_wb_clk_i;
 wire clknet_leaf_135_wb_clk_i;
 wire clknet_leaf_136_wb_clk_i;
 wire clknet_leaf_137_wb_clk_i;
 wire clknet_leaf_138_wb_clk_i;
 wire clknet_leaf_139_wb_clk_i;
 wire clknet_leaf_140_wb_clk_i;
 wire clknet_leaf_141_wb_clk_i;
 wire clknet_leaf_142_wb_clk_i;
 wire clknet_leaf_143_wb_clk_i;
 wire clknet_leaf_144_wb_clk_i;
 wire clknet_leaf_145_wb_clk_i;
 wire clknet_0_wb_clk_i;
 wire clknet_4_0_0_wb_clk_i;
 wire clknet_4_1_0_wb_clk_i;
 wire clknet_4_2_0_wb_clk_i;
 wire clknet_4_3_0_wb_clk_i;
 wire clknet_4_4_0_wb_clk_i;
 wire clknet_4_5_0_wb_clk_i;
 wire clknet_4_6_0_wb_clk_i;
 wire clknet_4_7_0_wb_clk_i;
 wire clknet_4_8_0_wb_clk_i;
 wire clknet_4_9_0_wb_clk_i;
 wire clknet_4_10_0_wb_clk_i;
 wire clknet_4_11_0_wb_clk_i;
 wire clknet_4_12_0_wb_clk_i;
 wire clknet_4_13_0_wb_clk_i;
 wire clknet_4_14_0_wb_clk_i;
 wire clknet_4_15_0_wb_clk_i;
 wire clknet_opt_1_0_wb_clk_i;

 gf180mcu_fd_sc_mcu7t5v0__inv_4 _3053_ (.I(net18),
    .ZN(_0674_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _3054_ (.I(_0674_),
    .Z(_0675_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3055_ (.I(_0675_),
    .Z(_0676_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _3056_ (.A1(\soc.spi_video_ram_1.state_counter[9] ),
    .A2(\soc.spi_video_ram_1.state_counter[8] ),
    .A3(\soc.spi_video_ram_1.state_counter[10] ),
    .ZN(_0677_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _3057_ (.A1(\soc.spi_video_ram_1.state_counter[5] ),
    .A2(\soc.spi_video_ram_1.state_counter[4] ),
    .A3(\soc.spi_video_ram_1.state_counter[7] ),
    .A4(\soc.spi_video_ram_1.state_counter[6] ),
    .ZN(_0678_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _3058_ (.A1(\soc.spi_video_ram_1.state_counter[1] ),
    .A2(\soc.spi_video_ram_1.state_counter[0] ),
    .A3(\soc.spi_video_ram_1.state_counter[3] ),
    .A4(\soc.spi_video_ram_1.state_counter[2] ),
    .ZN(_0679_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3059_ (.A1(_0677_),
    .A2(_0678_),
    .A3(_0679_),
    .ZN(_0680_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3060_ (.I(\soc.spi_video_ram_1.state_sram_clk_counter[1] ),
    .ZN(_0681_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _3061_ (.A1(\soc.spi_video_ram_1.state_sram_clk_counter[7] ),
    .A2(\soc.spi_video_ram_1.state_sram_clk_counter[6] ),
    .A3(\soc.spi_video_ram_1.state_sram_clk_counter[5] ),
    .A4(\soc.spi_video_ram_1.state_sram_clk_counter[4] ),
    .ZN(_0682_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3062_ (.A1(\soc.spi_video_ram_1.state_sram_clk_counter[3] ),
    .A2(\soc.spi_video_ram_1.state_sram_clk_counter[2] ),
    .ZN(_0683_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3063_ (.A1(_0682_),
    .A2(_0683_),
    .ZN(_0684_));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _3064_ (.A1(\soc.spi_video_ram_1.state_sram_clk_counter[8] ),
    .A2(\soc.spi_video_ram_1.state_sram_clk_counter[0] ),
    .A3(_0684_),
    .Z(_0685_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _3065_ (.A1(_0681_),
    .A2(_0685_),
    .ZN(_0686_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3066_ (.A1(_0680_),
    .A2(_0686_),
    .ZN(_0687_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3067_ (.A1(\soc.spi_video_ram_1.current_state[0] ),
    .A2(_0687_),
    .ZN(_0688_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3068_ (.A1(_0676_),
    .A2(_0688_),
    .ZN(_0003_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3069_ (.I(net18),
    .Z(_0689_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3070_ (.I(_0689_),
    .Z(_0690_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3071_ (.I(_0690_),
    .Z(_0691_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3072_ (.I(_0687_),
    .ZN(_0692_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3073_ (.I(\soc.spi_video_ram_1.write_fifo.write_pointer[0] ),
    .ZN(_0693_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 _3074_ (.I(\soc.spi_video_ram_1.write_fifo.write_pointer[1] ),
    .Z(_0694_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3075_ (.A1(\soc.spi_video_ram_1.write_fifo.read_pointer[1] ),
    .A2(_0694_),
    .Z(_0695_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3076_ (.A1(\soc.spi_video_ram_1.write_fifo.read_pointer[0] ),
    .A2(_0693_),
    .B(_0695_),
    .ZN(_0696_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3077_ (.I(\soc.spi_video_ram_1.write_fifo.read_pointer[0] ),
    .ZN(_0697_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _3078_ (.I(\soc.spi_video_ram_1.write_fifo.write_pointer[0] ),
    .Z(_0698_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3079_ (.A1(_0697_),
    .A2(_0698_),
    .ZN(_0699_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _3080_ (.I(\soc.spi_video_ram_1.write_fifo.write_pointer[2] ),
    .ZN(_0700_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3081_ (.A1(\soc.spi_video_ram_1.write_fifo.read_pointer[2] ),
    .A2(_0700_),
    .Z(_0701_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _3082_ (.A1(_0696_),
    .A2(_0699_),
    .A3(_0701_),
    .Z(_0702_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3083_ (.I(\soc.spi_video_ram_1.current_state[1] ),
    .Z(_0703_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _3084_ (.A1(_0703_),
    .A2(\soc.spi_video_ram_1.current_state[4] ),
    .Z(_0704_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _3085_ (.A1(\soc.spi_video_ram_1.current_state[3] ),
    .A2(\soc.spi_video_ram_1.current_state[0] ),
    .A3(_0704_),
    .ZN(_0705_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3086_ (.I(_0705_),
    .ZN(_0706_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3087_ (.A1(_0702_),
    .A2(_0706_),
    .B(\soc.spi_video_ram_1.initialized ),
    .ZN(_0707_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3088_ (.I(\soc.spi_video_ram_1.current_state[2] ),
    .ZN(_0708_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _3089_ (.A1(\soc.spi_video_ram_1.start_read ),
    .A2(_0702_),
    .B(_0707_),
    .C(_0708_),
    .ZN(_0709_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _3090_ (.I(_0703_),
    .ZN(_0710_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3091_ (.I(\soc.spi_video_ram_1.state_sram_clk_counter[2] ),
    .ZN(_0711_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _3092_ (.A1(\soc.spi_video_ram_1.state_sram_clk_counter[8] ),
    .A2(\soc.spi_video_ram_1.state_sram_clk_counter[1] ),
    .A3(\soc.spi_video_ram_1.state_sram_clk_counter[0] ),
    .ZN(_0712_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3093_ (.A1(\soc.spi_video_ram_1.state_sram_clk_counter[3] ),
    .A2(_0682_),
    .A3(_0712_),
    .ZN(_0713_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _3094_ (.A1(_0711_),
    .A2(_0713_),
    .Z(_0714_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _3095_ (.A1(\soc.spi_video_ram_1.state_sram_clk_counter[8] ),
    .A2(_0681_),
    .Z(_0715_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3096_ (.I(_0715_),
    .ZN(_0716_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3097_ (.A1(\soc.spi_video_ram_1.state_sram_clk_counter[3] ),
    .A2(_0711_),
    .A3(\soc.spi_video_ram_1.state_sram_clk_counter[0] ),
    .ZN(_0717_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _3098_ (.A1(\soc.spi_video_ram_1.state_sram_clk_counter[6] ),
    .A2(\soc.spi_video_ram_1.state_sram_clk_counter[5] ),
    .A3(\soc.spi_video_ram_1.state_sram_clk_counter[4] ),
    .A4(_0717_),
    .ZN(_0718_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _3099_ (.A1(\soc.spi_video_ram_1.state_sram_clk_counter[7] ),
    .A2(\soc.spi_video_ram_1.current_state[4] ),
    .A3(_0716_),
    .A4(_0718_),
    .ZN(_0719_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _3100_ (.I(\soc.spi_video_ram_1.current_state[3] ),
    .Z(_0720_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3101_ (.A1(\soc.spi_video_ram_1.state_sram_clk_counter[2] ),
    .A2(_0713_),
    .ZN(_0721_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3102_ (.A1(_0720_),
    .A2(_0721_),
    .ZN(_0722_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3103_ (.A1(_0710_),
    .A2(_0714_),
    .B(_0719_),
    .C(_0722_),
    .ZN(_0723_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _3104_ (.A1(\soc.spi_video_ram_1.current_state[0] ),
    .A2(_0692_),
    .B(_0709_),
    .C(_0723_),
    .ZN(_0724_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3105_ (.A1(_0691_),
    .A2(_0724_),
    .ZN(_0005_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _3106_ (.A1(\soc.spi_video_ram_1.state_sram_clk_counter[2] ),
    .A2(_0713_),
    .Z(_0725_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3107_ (.A1(\soc.spi_video_ram_1.current_state[3] ),
    .A2(_0725_),
    .ZN(_0726_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3108_ (.I(\soc.spi_video_ram_1.initialized ),
    .ZN(_0727_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3109_ (.A1(_0727_),
    .A2(\soc.spi_video_ram_1.current_state[2] ),
    .ZN(_0728_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3110_ (.A1(_0726_),
    .A2(_0728_),
    .B(_0691_),
    .ZN(_0006_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3111_ (.I(\soc.spi_video_ram_1.current_state[4] ),
    .Z(_0729_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3112_ (.A1(\soc.spi_video_ram_1.state_sram_clk_counter[5] ),
    .A2(\soc.spi_video_ram_1.state_sram_clk_counter[4] ),
    .ZN(_0730_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3113_ (.A1(\soc.spi_video_ram_1.state_sram_clk_counter[7] ),
    .A2(_0730_),
    .ZN(_0731_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _3114_ (.A1(\soc.spi_video_ram_1.state_sram_clk_counter[6] ),
    .A2(_0715_),
    .A3(_0717_),
    .A4(_0731_),
    .Z(_0732_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3115_ (.A1(_0729_),
    .A2(_0732_),
    .ZN(_0733_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _3116_ (.A1(\soc.spi_video_ram_1.initialized ),
    .A2(\soc.spi_video_ram_1.start_read ),
    .A3(\soc.spi_video_ram_1.current_state[2] ),
    .A4(_0702_),
    .ZN(_0734_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3117_ (.A1(_0733_),
    .A2(_0734_),
    .B(_0691_),
    .ZN(_0007_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3118_ (.A1(_0703_),
    .A2(_0714_),
    .ZN(_0735_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _3119_ (.A1(_0708_),
    .A2(_0702_),
    .A3(_0706_),
    .ZN(_0736_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3120_ (.I(_0736_),
    .Z(_0008_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3121_ (.A1(\soc.spi_video_ram_1.initialized ),
    .A2(_0008_),
    .ZN(_0737_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3122_ (.A1(_0735_),
    .A2(_0737_),
    .B(_0691_),
    .ZN(_0004_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3123_ (.A1(_0694_),
    .A2(\soc.spi_video_ram_1.write_fifo.write_pointer[0] ),
    .ZN(_0738_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3124_ (.A1(_0701_),
    .A2(_0738_),
    .Z(_0739_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _3125_ (.A1(_0695_),
    .A2(_0699_),
    .B(_0739_),
    .C(_0696_),
    .ZN(_0740_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _3126_ (.A1(\soc.rom_encoder_0.write_enable ),
    .A2(net18),
    .A3(net13),
    .A4(net37),
    .Z(_0741_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3127_ (.A1(\soc.ram_encoder_0.initialized ),
    .A2(\soc.rom_encoder_0.initialized ),
    .A3(\soc.spi_video_ram_1.initialized ),
    .ZN(_0742_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _3128_ (.A1(\soc.hack_wait_clocks[1] ),
    .A2(\soc.hack_wait_clocks[0] ),
    .A3(_0741_),
    .A4(_0742_),
    .Z(_0743_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3129_ (.A1(\soc.cpu.instruction[15] ),
    .A2(\soc.cpu.instruction[3] ),
    .ZN(_0744_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3130_ (.I(\soc.cpu.AReg.data[13] ),
    .ZN(_0745_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _3131_ (.A1(net87),
    .A2(\soc.hack_clk_strobe ),
    .A3(\soc.cpu.AReg.data[14] ),
    .A4(_0745_),
    .ZN(_0746_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _3132_ (.A1(_0740_),
    .A2(_0743_),
    .A3(_0744_),
    .A4(_0746_),
    .ZN(_0747_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 _3133_ (.I(_0747_),
    .Z(_0748_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3134_ (.I(_0748_),
    .Z(_0009_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _3135_ (.I(\soc.spi_video_ram_1.buffer_index[4] ),
    .ZN(_0749_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _3136_ (.I(\soc.spi_video_ram_1.buffer_index[0] ),
    .Z(_0750_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3137_ (.A1(_0750_),
    .A2(\soc.spi_video_ram_1.buffer_index[1] ),
    .ZN(_0751_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3138_ (.I(\soc.spi_video_ram_1.buffer_index[3] ),
    .Z(_0752_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _3139_ (.A1(\soc.spi_video_ram_1.buffer_index[2] ),
    .A2(_0752_),
    .ZN(_0753_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3140_ (.A1(\soc.spi_video_ram_1.buffer_index[4] ),
    .A2(_0753_),
    .Z(_0754_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3141_ (.A1(_0751_),
    .A2(_0754_),
    .ZN(_0755_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3142_ (.A1(_0749_),
    .A2(_0751_),
    .B(_0755_),
    .ZN(_0756_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _3143_ (.I(_0750_),
    .Z(_0757_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3144_ (.I(\soc.spi_video_ram_1.buffer_index[1] ),
    .Z(_0758_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3145_ (.I(\soc.spi_video_ram_1.buffer_index[2] ),
    .Z(_0759_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _3146_ (.A1(_0758_),
    .A2(_0759_),
    .Z(_0760_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _3147_ (.A1(_0750_),
    .A2(\soc.spi_video_ram_1.buffer_index[1] ),
    .B(_0759_),
    .ZN(_0761_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _3148_ (.A1(_0757_),
    .A2(_0760_),
    .B(_0761_),
    .ZN(_0762_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3149_ (.A1(\soc.spi_video_ram_1.buffer_index[0] ),
    .A2(\soc.spi_video_ram_1.buffer_index[1] ),
    .ZN(_0763_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _3150_ (.A1(_0750_),
    .A2(\soc.spi_video_ram_1.buffer_index[1] ),
    .Z(_0764_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3151_ (.A1(_0751_),
    .A2(_0764_),
    .Z(_0765_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3152_ (.I0(\soc.spi_video_ram_1.output_buffer[3] ),
    .I1(\soc.spi_video_ram_1.output_buffer[2] ),
    .S(_0750_),
    .Z(_0766_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3153_ (.A1(\soc.spi_video_ram_1.output_buffer[1] ),
    .A2(_0763_),
    .B1(_0765_),
    .B2(_0766_),
    .ZN(_0767_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3154_ (.I(_0767_),
    .ZN(_0768_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3155_ (.I(\soc.spi_video_ram_1.buffer_index[5] ),
    .ZN(_0769_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3156_ (.A1(_0749_),
    .A2(_0769_),
    .A3(_0753_),
    .ZN(_0770_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3157_ (.A1(\soc.spi_video_ram_1.buffer_index[1] ),
    .A2(_0770_),
    .ZN(_0771_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _3158_ (.A1(_0750_),
    .A2(_0771_),
    .ZN(_0772_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3159_ (.A1(_0757_),
    .A2(\soc.spi_video_ram_1.output_buffer[6] ),
    .B1(_0772_),
    .B2(\soc.spi_video_ram_1.output_buffer[7] ),
    .ZN(_0773_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3160_ (.A1(_0765_),
    .A2(_0773_),
    .B(_0762_),
    .ZN(_0774_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3161_ (.A1(_0751_),
    .A2(_0764_),
    .ZN(_0775_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3162_ (.I(_0750_),
    .Z(_0776_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3163_ (.A1(_0776_),
    .A2(\soc.spi_video_ram_1.output_buffer[4] ),
    .B1(_0772_),
    .B2(\soc.spi_video_ram_1.output_buffer[5] ),
    .ZN(_0777_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3164_ (.A1(_0775_),
    .A2(_0777_),
    .ZN(_0778_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3165_ (.I(_0761_),
    .ZN(_0779_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3166_ (.A1(_0752_),
    .A2(_0779_),
    .Z(_0780_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3167_ (.I(_0780_),
    .ZN(_0781_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _3168_ (.A1(_0762_),
    .A2(_0768_),
    .B1(_0774_),
    .B2(_0778_),
    .C(_0781_),
    .ZN(_0782_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 _3169_ (.I(_0750_),
    .Z(_0783_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3170_ (.I0(\soc.spi_video_ram_1.output_buffer[11] ),
    .I1(\soc.spi_video_ram_1.output_buffer[10] ),
    .S(_0783_),
    .Z(_0784_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3171_ (.I0(\soc.spi_video_ram_1.output_buffer[9] ),
    .I1(\soc.spi_video_ram_1.output_buffer[8] ),
    .S(_0783_),
    .Z(_0785_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3172_ (.I0(_0784_),
    .I1(_0785_),
    .S(_0775_),
    .Z(_0786_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3173_ (.A1(_0776_),
    .A2(\soc.spi_video_ram_1.output_buffer[12] ),
    .B1(_0772_),
    .B2(\soc.spi_video_ram_1.output_buffer[13] ),
    .ZN(_0787_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3174_ (.A1(_0783_),
    .A2(\soc.spi_video_ram_1.output_buffer[14] ),
    .ZN(_0788_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3175_ (.A1(\soc.spi_video_ram_1.output_buffer[15] ),
    .A2(_0770_),
    .ZN(_0789_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _3176_ (.A1(_0771_),
    .A2(_0788_),
    .B1(_0789_),
    .B2(_0757_),
    .ZN(_0790_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3177_ (.A1(_0775_),
    .A2(_0790_),
    .ZN(_0791_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _3178_ (.A1(_0775_),
    .A2(_0787_),
    .B(_0791_),
    .C(_0762_),
    .ZN(_0792_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _3179_ (.A1(_0762_),
    .A2(_0786_),
    .B(_0792_),
    .C(_0780_),
    .ZN(_0793_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3180_ (.A1(_0776_),
    .A2(\soc.spi_video_ram_1.output_buffer[22] ),
    .B1(_0772_),
    .B2(\soc.spi_video_ram_1.output_buffer[23] ),
    .ZN(_0794_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3181_ (.A1(_0775_),
    .A2(_0794_),
    .ZN(_0795_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3182_ (.A1(_0776_),
    .A2(\soc.spi_video_ram_1.output_buffer[20] ),
    .B1(_0772_),
    .B2(\soc.spi_video_ram_1.output_buffer[21] ),
    .ZN(_0796_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3183_ (.A1(_0765_),
    .A2(_0796_),
    .ZN(_0797_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _3184_ (.A1(_0762_),
    .A2(_0795_),
    .A3(_0797_),
    .ZN(_0798_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3185_ (.I(\soc.spi_video_ram_1.output_buffer[17] ),
    .ZN(_0799_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3186_ (.I(\soc.spi_video_ram_1.output_buffer[19] ),
    .ZN(_0800_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3187_ (.I(\soc.spi_video_ram_1.output_buffer[18] ),
    .ZN(_0801_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3188_ (.I(\soc.spi_video_ram_1.output_buffer[16] ),
    .ZN(_0802_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3189_ (.I0(_0799_),
    .I1(_0800_),
    .I2(_0801_),
    .I3(_0802_),
    .S0(_0758_),
    .S1(_0776_),
    .Z(_0803_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3190_ (.A1(_0762_),
    .A2(_0803_),
    .ZN(_0804_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3191_ (.A1(\soc.spi_video_ram_1.buffer_index[4] ),
    .A2(_0780_),
    .A3(_0804_),
    .ZN(_0805_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _3192_ (.A1(_0756_),
    .A2(_0782_),
    .A3(_0793_),
    .B1(_0798_),
    .B2(_0805_),
    .ZN(_0806_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3193_ (.A1(_0720_),
    .A2(\soc.spi_video_ram_1.buffer_index[5] ),
    .ZN(_0807_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _3194_ (.A1(_0758_),
    .A2(_0759_),
    .ZN(_0808_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3195_ (.I0(\soc.spi_video_ram_1.output_buffer[8] ),
    .I1(\soc.spi_video_ram_1.output_buffer[9] ),
    .S(_0783_),
    .Z(_0809_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3196_ (.I(_0759_),
    .ZN(_0810_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3197_ (.A1(_0758_),
    .A2(_0810_),
    .Z(_0811_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3198_ (.I0(\soc.spi_video_ram_1.output_buffer[10] ),
    .I1(\soc.spi_video_ram_1.output_buffer[11] ),
    .S(_0757_),
    .Z(_0812_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3199_ (.A1(_0808_),
    .A2(_0809_),
    .B1(_0811_),
    .B2(_0812_),
    .ZN(_0813_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3200_ (.I0(\soc.spi_video_ram_1.output_buffer[14] ),
    .I1(\soc.spi_video_ram_1.output_buffer[15] ),
    .S(_0783_),
    .Z(_0814_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _3201_ (.A1(_0758_),
    .A2(_0810_),
    .ZN(_0815_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3202_ (.I0(\soc.spi_video_ram_1.output_buffer[12] ),
    .I1(\soc.spi_video_ram_1.output_buffer[13] ),
    .S(_0783_),
    .Z(_0816_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3203_ (.A1(_0760_),
    .A2(_0814_),
    .B1(_0815_),
    .B2(_0816_),
    .ZN(_0817_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3204_ (.A1(_0813_),
    .A2(_0817_),
    .ZN(_0818_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3205_ (.A1(_0752_),
    .A2(_0818_),
    .ZN(_0819_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3206_ (.I(\soc.spi_video_ram_1.output_buffer[22] ),
    .ZN(_0820_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3207_ (.A1(_0757_),
    .A2(\soc.spi_video_ram_1.output_buffer[23] ),
    .ZN(_0821_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3208_ (.A1(_0776_),
    .A2(_0820_),
    .B(_0821_),
    .ZN(_0822_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3209_ (.A1(_0760_),
    .A2(_0822_),
    .ZN(_0823_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3210_ (.A1(_0783_),
    .A2(\soc.spi_video_ram_1.output_buffer[17] ),
    .ZN(_0824_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3211_ (.A1(_0757_),
    .A2(_0802_),
    .B(_0824_),
    .ZN(_0825_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3212_ (.A1(_0783_),
    .A2(\soc.spi_video_ram_1.output_buffer[19] ),
    .ZN(_0826_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3213_ (.A1(_0757_),
    .A2(_0801_),
    .B(_0826_),
    .ZN(_0827_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3214_ (.I(\soc.spi_video_ram_1.output_buffer[20] ),
    .ZN(_0828_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3215_ (.A1(_0783_),
    .A2(\soc.spi_video_ram_1.output_buffer[21] ),
    .ZN(_0829_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3216_ (.A1(_0757_),
    .A2(_0828_),
    .B(_0829_),
    .ZN(_0830_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _3217_ (.A1(_0808_),
    .A2(_0825_),
    .B1(_0827_),
    .B2(_0811_),
    .C1(_0815_),
    .C2(_0830_),
    .ZN(_0831_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3218_ (.A1(\soc.spi_video_ram_1.buffer_index[4] ),
    .A2(_0823_),
    .A3(_0831_),
    .ZN(_0832_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3219_ (.I(\soc.spi_video_ram_1.output_buffer[4] ),
    .ZN(_0833_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3220_ (.A1(_0783_),
    .A2(\soc.spi_video_ram_1.output_buffer[5] ),
    .ZN(_0834_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3221_ (.A1(_0757_),
    .A2(_0833_),
    .B(_0834_),
    .C(_0759_),
    .ZN(_0835_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3222_ (.I(_0835_),
    .ZN(_0836_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3223_ (.A1(_0776_),
    .A2(\soc.spi_video_ram_1.output_buffer[1] ),
    .B(_0759_),
    .ZN(_0837_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3224_ (.I0(\soc.spi_video_ram_1.output_buffer[6] ),
    .I1(\soc.spi_video_ram_1.output_buffer[7] ),
    .S(_0750_),
    .Z(_0838_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3225_ (.I0(\soc.spi_video_ram_1.output_buffer[2] ),
    .I1(\soc.spi_video_ram_1.output_buffer[3] ),
    .S(_0750_),
    .Z(_0839_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _3226_ (.A1(_0760_),
    .A2(_0838_),
    .B1(_0839_),
    .B2(_0811_),
    .C(\soc.spi_video_ram_1.buffer_index[4] ),
    .ZN(_0840_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _3227_ (.A1(_0758_),
    .A2(_0836_),
    .A3(_0837_),
    .B(_0840_),
    .ZN(_0841_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3228_ (.A1(_0832_),
    .A2(_0841_),
    .ZN(_0842_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _3229_ (.A1(\soc.spi_video_ram_1.buffer_index[4] ),
    .A2(_0819_),
    .B1(_0842_),
    .B2(_0752_),
    .ZN(_0843_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3230_ (.A1(_0806_),
    .A2(_0807_),
    .B1(_0843_),
    .B2(_0720_),
    .ZN(_0844_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3231_ (.I(_0844_),
    .ZN(net70));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3232_ (.I(\soc.cpu.instruction[15] ),
    .Z(_0845_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _3233_ (.I(_0845_),
    .Z(_0846_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3234_ (.I(\soc.cpu.DMuxJMP.sel[0] ),
    .ZN(_0847_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3235_ (.A1(_0845_),
    .A2(\soc.cpu.instruction[5] ),
    .ZN(_0848_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _3236_ (.I(\soc.cpu.ALU.nx ),
    .Z(_0849_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _3237_ (.I(\soc.cpu.ALU.zx ),
    .ZN(_0850_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3238_ (.A1(_0850_),
    .A2(\soc.cpu.ALU.x[0] ),
    .ZN(_0851_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3239_ (.A1(_0849_),
    .A2(_0851_),
    .Z(_0852_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _3240_ (.I(\soc.cpu.ALU.ny ),
    .Z(_0853_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _3241_ (.I(\soc.cpu.instruction[12] ),
    .ZN(_0854_));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 _3242_ (.I(\soc.cpu.AReg.data[0] ),
    .ZN(_0855_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _3243_ (.A1(\soc.cpu.AReg.data[4] ),
    .A2(\soc.cpu.AReg.data[7] ),
    .A3(\soc.cpu.AReg.data[6] ),
    .ZN(_0856_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _3244_ (.A1(\soc.cpu.AReg.data[11] ),
    .A2(\soc.cpu.AReg.data[10] ),
    .A3(\soc.cpu.AReg.data[12] ),
    .A4(\soc.cpu.AReg.data[5] ),
    .ZN(_0857_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3245_ (.A1(\soc.cpu.AReg.data[14] ),
    .A2(\soc.cpu.AReg.data[13] ),
    .Z(_0858_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3246_ (.A1(\soc.cpu.AReg.data[9] ),
    .A2(\soc.cpu.AReg.data[8] ),
    .ZN(_0859_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _3247_ (.A1(_0856_),
    .A2(_0857_),
    .A3(_0858_),
    .A4(_0859_),
    .Z(_0860_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3248_ (.A1(\soc.cpu.AReg.data[3] ),
    .A2(\soc.cpu.AReg.data[2] ),
    .ZN(_0861_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3249_ (.A1(\soc.cpu.AReg.data[1] ),
    .A2(_0861_),
    .Z(_0862_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _3250_ (.A1(net77),
    .A2(_0855_),
    .A3(_0860_),
    .A4(_0862_),
    .ZN(_0863_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _3251_ (.A1(_0856_),
    .A2(_0857_),
    .A3(_0858_),
    .A4(_0859_),
    .ZN(_0864_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _3252_ (.A1(\soc.cpu.AReg.data[3] ),
    .A2(\soc.cpu.AReg.data[2] ),
    .A3(\soc.cpu.AReg.data[1] ),
    .ZN(_0865_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _3253_ (.I(_0865_),
    .ZN(_0866_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _3254_ (.A1(_0855_),
    .A2(_0864_),
    .A3(_0866_),
    .ZN(_0867_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _3255_ (.A1(\soc.cpu.AReg.data[0] ),
    .A2(_0864_),
    .A3(_0866_),
    .ZN(_0868_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _3256_ (.A1(\soc.cpu.AReg.data[14] ),
    .A2(\soc.cpu.AReg.data[13] ),
    .ZN(_0869_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3257_ (.A1(\soc.ram_data_out[0] ),
    .A2(_0869_),
    .ZN(_0870_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3258_ (.A1(\soc.cpu.instruction[12] ),
    .A2(_0870_),
    .ZN(_0871_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _3259_ (.A1(\soc.gpio_i_stored[0] ),
    .A2(_0867_),
    .B1(_0868_),
    .B2(net29),
    .C(_0871_),
    .ZN(_0872_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _3260_ (.A1(_0854_),
    .A2(_0855_),
    .B1(_0863_),
    .B2(_0872_),
    .C(\soc.cpu.ALU.zy ),
    .ZN(_0873_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3261_ (.A1(_0853_),
    .A2(_0873_),
    .ZN(_0874_));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 _3262_ (.I(\soc.cpu.ALU.f ),
    .ZN(_0875_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3263_ (.A1(_0852_),
    .A2(_0874_),
    .B(_0875_),
    .ZN(_0876_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3264_ (.A1(_0852_),
    .A2(_0874_),
    .ZN(_0877_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _3265_ (.A1(\soc.cpu.ALU.no ),
    .A2(_0876_),
    .A3(_0877_),
    .ZN(_0878_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3266_ (.I(\soc.cpu.instruction[5] ),
    .ZN(_0879_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3267_ (.A1(\soc.cpu.instruction[15] ),
    .A2(_0879_),
    .ZN(_0880_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3268_ (.I(_0880_),
    .Z(_0881_));
 gf180mcu_fd_sc_mcu7t5v0__oai222_2 _3269_ (.A1(_0846_),
    .A2(_0847_),
    .B1(_0848_),
    .B2(_0878_),
    .C1(_0881_),
    .C2(_0855_),
    .ZN(\soc.cpu.PC.in[0] ));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3270_ (.A1(\soc.cpu.instruction[15] ),
    .A2(\soc.cpu.instruction[5] ),
    .Z(_0882_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3271_ (.I(_0882_),
    .Z(_0883_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3272_ (.I(_0883_),
    .Z(_0884_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3273_ (.A1(_0850_),
    .A2(\soc.cpu.ALU.x[1] ),
    .ZN(_0885_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3274_ (.A1(_0849_),
    .A2(_0885_),
    .Z(_0886_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _3275_ (.I(\soc.cpu.instruction[12] ),
    .Z(_0887_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3276_ (.A1(\soc.ram_data_out[1] ),
    .A2(_0869_),
    .ZN(_0888_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3277_ (.A1(_0887_),
    .A2(_0888_),
    .ZN(_0889_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3278_ (.I(net38),
    .ZN(_0890_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _3279_ (.A1(net78),
    .A2(_0855_),
    .A3(_0860_),
    .A4(_0862_),
    .ZN(_0891_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3280_ (.A1(\soc.gpio_i_stored[1] ),
    .A2(_0855_),
    .B(_0860_),
    .C(_0865_),
    .ZN(_0892_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _3281_ (.A1(_0890_),
    .A2(_0868_),
    .B1(_0891_),
    .B2(_0892_),
    .C(_0869_),
    .ZN(_0893_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _3282_ (.I(\soc.cpu.ALU.zy ),
    .ZN(_0894_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _3283_ (.A1(_0887_),
    .A2(\soc.cpu.AReg.data[1] ),
    .B1(_0889_),
    .B2(_0893_),
    .C(_0894_),
    .ZN(_0895_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _3284_ (.A1(_0853_),
    .A2(_0886_),
    .A3(_0895_),
    .ZN(_0896_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3285_ (.A1(_0877_),
    .A2(_0896_),
    .Z(_0897_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3286_ (.A1(\soc.cpu.ALU.f ),
    .A2(_0897_),
    .ZN(_0898_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3287_ (.A1(_0853_),
    .A2(_0895_),
    .Z(_0899_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3288_ (.A1(_0886_),
    .A2(_0899_),
    .B(_0875_),
    .ZN(_0900_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3289_ (.A1(_0898_),
    .A2(_0900_),
    .Z(_0901_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _3290_ (.A1(\soc.cpu.ALU.no ),
    .A2(_0901_),
    .ZN(_0902_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _3291_ (.A1(_0846_),
    .A2(\soc.cpu.DMuxJMP.sel[1] ),
    .B1(\soc.cpu.AReg.data[1] ),
    .B2(_0881_),
    .ZN(_0903_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3292_ (.A1(_0884_),
    .A2(_0902_),
    .B(_0903_),
    .ZN(\soc.cpu.PC.in[1] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3293_ (.I(_0850_),
    .Z(_0904_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3294_ (.A1(_0904_),
    .A2(\soc.cpu.ALU.x[2] ),
    .ZN(_0905_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3295_ (.A1(_0849_),
    .A2(_0905_),
    .ZN(_0906_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3296_ (.I(_0854_),
    .Z(_0907_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3297_ (.I(\soc.cpu.AReg.data[2] ),
    .ZN(_0908_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3298_ (.A1(\soc.ram_data_out[2] ),
    .A2(_0869_),
    .B(_0854_),
    .ZN(_0909_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _3299_ (.A1(net79),
    .A2(_0855_),
    .A3(_0860_),
    .A4(_0862_),
    .Z(_0910_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _3300_ (.A1(\soc.gpio_i_stored[2] ),
    .A2(\soc.cpu.AReg.data[0] ),
    .A3(_0860_),
    .A4(_0865_),
    .Z(_0911_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _3301_ (.A1(\soc.cpu.AReg.data[0] ),
    .A2(net39),
    .A3(_0864_),
    .A4(_0866_),
    .Z(_0912_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _3302_ (.A1(_0868_),
    .A2(_0910_),
    .A3(_0911_),
    .B(_0912_),
    .ZN(_0913_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _3303_ (.A1(_0907_),
    .A2(_0908_),
    .B1(_0909_),
    .B2(_0913_),
    .C(\soc.cpu.ALU.zy ),
    .ZN(_0914_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3304_ (.A1(_0853_),
    .A2(_0914_),
    .Z(_0915_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3305_ (.A1(_0906_),
    .A2(_0915_),
    .Z(_0916_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _3306_ (.A1(_0852_),
    .A2(_0874_),
    .A3(_0896_),
    .B1(_0899_),
    .B2(_0886_),
    .ZN(_0917_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _3307_ (.A1(_0917_),
    .A2(_0906_),
    .A3(_0915_),
    .Z(_0918_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3308_ (.I0(_0916_),
    .I1(_0918_),
    .S(\soc.cpu.ALU.f ),
    .Z(_0919_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _3309_ (.A1(\soc.cpu.ALU.no ),
    .A2(_0919_),
    .ZN(_0920_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _3310_ (.A1(_0846_),
    .A2(\soc.cpu.DMuxJMP.sel[2] ),
    .B1(\soc.cpu.AReg.data[2] ),
    .B2(_0881_),
    .ZN(_0921_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3311_ (.A1(_0884_),
    .A2(_0920_),
    .B(_0921_),
    .ZN(\soc.cpu.PC.in[2] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _3312_ (.I(\soc.cpu.ALU.no ),
    .Z(_0922_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _3313_ (.I(_0849_),
    .Z(_0923_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3314_ (.A1(_0904_),
    .A2(\soc.cpu.ALU.x[3] ),
    .ZN(_0924_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3315_ (.A1(_0923_),
    .A2(_0924_),
    .ZN(_0925_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _3316_ (.I(_0853_),
    .Z(_0926_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3317_ (.A1(\soc.ram_data_out[3] ),
    .A2(_0869_),
    .ZN(_0927_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3318_ (.A1(_0887_),
    .A2(_0927_),
    .ZN(_0928_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3319_ (.I(net40),
    .ZN(_0929_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3320_ (.A1(\soc.cpu.AReg.data[1] ),
    .A2(_0861_),
    .ZN(_0930_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _3321_ (.A1(\soc.cpu.AReg.data[0] ),
    .A2(_0864_),
    .A3(_0930_),
    .ZN(_0931_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _3322_ (.A1(net80),
    .A2(_0931_),
    .B1(_0867_),
    .B2(\soc.gpio_i_stored[3] ),
    .C(_0868_),
    .ZN(_0932_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3323_ (.A1(_0929_),
    .A2(_0868_),
    .B(_0932_),
    .ZN(_0933_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _3324_ (.A1(_0887_),
    .A2(\soc.cpu.AReg.data[3] ),
    .B1(_0928_),
    .B2(_0933_),
    .C(_0894_),
    .ZN(_0934_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3325_ (.A1(_0926_),
    .A2(_0934_),
    .ZN(_0935_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _3326_ (.A1(_0906_),
    .A2(_0915_),
    .Z(_0936_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _3327_ (.A1(_0917_),
    .A2(_0936_),
    .B(_0916_),
    .ZN(_0937_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _3328_ (.A1(_0925_),
    .A2(_0935_),
    .A3(_0937_),
    .ZN(_0938_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3329_ (.A1(_0925_),
    .A2(_0935_),
    .ZN(_0939_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3330_ (.A1(_0875_),
    .A2(_0939_),
    .ZN(_0940_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3331_ (.A1(_0875_),
    .A2(_0938_),
    .B(_0940_),
    .ZN(_0941_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _3332_ (.A1(_0922_),
    .A2(_0941_),
    .Z(_0942_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _3333_ (.A1(_0845_),
    .A2(\soc.cpu.instruction[3] ),
    .B1(\soc.cpu.AReg.data[3] ),
    .B2(_0881_),
    .ZN(_0943_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3334_ (.A1(_0884_),
    .A2(_0942_),
    .B(_0943_),
    .ZN(\soc.cpu.PC.in[3] ));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3335_ (.A1(_0925_),
    .A2(_0935_),
    .ZN(_0944_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _3336_ (.A1(_0937_),
    .A2(_0944_),
    .B(_0939_),
    .ZN(_0945_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3337_ (.A1(_0850_),
    .A2(\soc.cpu.ALU.x[4] ),
    .ZN(_0946_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3338_ (.A1(_0849_),
    .A2(_0946_),
    .ZN(_0947_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _3339_ (.A1(\soc.ram_data_out[4] ),
    .A2(_0869_),
    .B1(_0868_),
    .B2(net41),
    .C(_0854_),
    .ZN(_0948_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3340_ (.A1(_0887_),
    .A2(\soc.cpu.AReg.data[4] ),
    .B(_0894_),
    .ZN(_0949_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3341_ (.A1(_0948_),
    .A2(_0949_),
    .ZN(_0950_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3342_ (.A1(_0853_),
    .A2(_0950_),
    .Z(_0951_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3343_ (.A1(_0947_),
    .A2(_0951_),
    .Z(_0952_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3344_ (.A1(_0945_),
    .A2(_0952_),
    .Z(_0953_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3345_ (.I(\soc.cpu.ALU.f ),
    .Z(_0954_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3346_ (.A1(_0947_),
    .A2(_0951_),
    .Z(_0955_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _3347_ (.A1(_0954_),
    .A2(_0955_),
    .Z(_0956_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3348_ (.A1(_0875_),
    .A2(_0953_),
    .B(_0956_),
    .ZN(_0957_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3349_ (.A1(_0922_),
    .A2(_0957_),
    .Z(_0958_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _3350_ (.A1(_0846_),
    .A2(\soc.cpu.instruction[4] ),
    .B1(\soc.cpu.AReg.data[4] ),
    .B2(_0881_),
    .ZN(_0959_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3351_ (.A1(_0884_),
    .A2(_0958_),
    .B(_0959_),
    .ZN(\soc.cpu.PC.in[4] ));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _3352_ (.A1(_0945_),
    .A2(_0952_),
    .B(_0955_),
    .C(_0875_),
    .ZN(_0960_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3353_ (.A1(_0904_),
    .A2(\soc.cpu.ALU.x[5] ),
    .ZN(_0961_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3354_ (.A1(_0923_),
    .A2(_0961_),
    .ZN(_0962_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _3355_ (.A1(\soc.ram_data_out[5] ),
    .A2(_0869_),
    .B1(_0868_),
    .B2(net42),
    .C(_0907_),
    .ZN(_0963_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3356_ (.A1(_0887_),
    .A2(\soc.cpu.AReg.data[5] ),
    .B(_0894_),
    .ZN(_0964_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3357_ (.A1(_0963_),
    .A2(_0964_),
    .ZN(_0965_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3358_ (.A1(_0926_),
    .A2(_0965_),
    .Z(_0966_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3359_ (.A1(_0962_),
    .A2(_0966_),
    .ZN(_0967_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3360_ (.A1(_0962_),
    .A2(_0966_),
    .Z(_0968_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3361_ (.A1(_0954_),
    .A2(_0967_),
    .B(_0968_),
    .ZN(_0969_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _3362_ (.A1(_0922_),
    .A2(_0960_),
    .A3(_0969_),
    .Z(_0970_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3363_ (.A1(_0846_),
    .A2(\soc.cpu.AReg.data[5] ),
    .ZN(_0971_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3364_ (.A1(_0884_),
    .A2(_0970_),
    .B1(_0971_),
    .B2(_0879_),
    .ZN(\soc.cpu.PC.in[5] ));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3365_ (.I(_0875_),
    .Z(_0972_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3366_ (.A1(_0850_),
    .A2(\soc.cpu.ALU.x[6] ),
    .ZN(_0973_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3367_ (.A1(_0849_),
    .A2(_0973_),
    .ZN(_0974_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _3368_ (.A1(\soc.ram_data_out[6] ),
    .A2(_0869_),
    .B1(_0868_),
    .B2(net43),
    .C(_0854_),
    .ZN(_0975_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3369_ (.A1(_0887_),
    .A2(\soc.cpu.AReg.data[6] ),
    .B(_0894_),
    .ZN(_0976_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3370_ (.A1(_0975_),
    .A2(_0976_),
    .ZN(_0977_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3371_ (.A1(_0853_),
    .A2(_0977_),
    .Z(_0978_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3372_ (.A1(_0974_),
    .A2(_0978_),
    .ZN(_0979_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3373_ (.I(_0952_),
    .ZN(_0980_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _3374_ (.A1(_0980_),
    .A2(_0968_),
    .A3(_0967_),
    .ZN(_0981_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3375_ (.A1(_0947_),
    .A2(_0951_),
    .B1(_0962_),
    .B2(_0966_),
    .ZN(_0982_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3376_ (.A1(_0967_),
    .A2(_0982_),
    .ZN(_0983_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3377_ (.A1(_0945_),
    .A2(_0981_),
    .B(_0983_),
    .ZN(_0984_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3378_ (.A1(_0979_),
    .A2(_0984_),
    .Z(_0985_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3379_ (.A1(_0974_),
    .A2(_0978_),
    .ZN(_0986_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3380_ (.A1(_0875_),
    .A2(_0986_),
    .ZN(_0987_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3381_ (.A1(_0972_),
    .A2(_0985_),
    .B(_0987_),
    .ZN(_0988_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3382_ (.A1(_0922_),
    .A2(_0988_),
    .Z(_0989_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _3383_ (.I(_0922_),
    .Z(_0990_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _3384_ (.A1(_0846_),
    .A2(_0990_),
    .B1(\soc.cpu.AReg.data[6] ),
    .B2(_0881_),
    .ZN(_0991_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3385_ (.A1(_0884_),
    .A2(_0989_),
    .B(_0991_),
    .ZN(\soc.cpu.PC.in[6] ));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3386_ (.A1(_0979_),
    .A2(_0984_),
    .B(\soc.cpu.ALU.f ),
    .C(_0986_),
    .ZN(_0992_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3387_ (.A1(_0904_),
    .A2(\soc.cpu.ALU.x[7] ),
    .ZN(_0993_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3388_ (.A1(_0849_),
    .A2(_0993_),
    .ZN(_0994_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _3389_ (.A1(\soc.ram_data_out[7] ),
    .A2(_0869_),
    .B1(_0868_),
    .B2(net44),
    .C(_0854_),
    .ZN(_0995_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3390_ (.A1(_0887_),
    .A2(\soc.cpu.AReg.data[7] ),
    .B(_0894_),
    .ZN(_0996_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3391_ (.A1(_0995_),
    .A2(_0996_),
    .ZN(_0997_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3392_ (.A1(_0853_),
    .A2(_0997_),
    .Z(_0998_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3393_ (.A1(_0994_),
    .A2(_0998_),
    .ZN(_0999_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3394_ (.A1(_0994_),
    .A2(_0998_),
    .Z(_1000_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3395_ (.A1(_0954_),
    .A2(_0999_),
    .B(_1000_),
    .ZN(_1001_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_2 _3396_ (.A1(_0922_),
    .A2(_0992_),
    .A3(_1001_),
    .ZN(_1002_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _3397_ (.A1(_0845_),
    .A2(_0954_),
    .B1(\soc.cpu.AReg.data[7] ),
    .B2(_0881_),
    .ZN(_1003_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3398_ (.A1(_0884_),
    .A2(_1002_),
    .B(_1003_),
    .ZN(\soc.cpu.PC.in[7] ));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _3399_ (.A1(_0979_),
    .A2(_1000_),
    .A3(_0999_),
    .ZN(_1004_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _3400_ (.A1(_0945_),
    .A2(_0981_),
    .A3(_1004_),
    .Z(_1005_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3401_ (.A1(_0983_),
    .A2(_1004_),
    .Z(_1006_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3402_ (.A1(_0986_),
    .A2(_0999_),
    .ZN(_1007_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _3403_ (.A1(_1000_),
    .A2(_1006_),
    .A3(_1007_),
    .Z(_1008_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3404_ (.A1(_0850_),
    .A2(\soc.cpu.ALU.x[8] ),
    .ZN(_1009_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3405_ (.A1(_0849_),
    .A2(_1009_),
    .ZN(_1010_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3406_ (.I(\soc.cpu.ALU.zy ),
    .Z(_1011_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _3407_ (.A1(_0854_),
    .A2(_0858_),
    .ZN(_1012_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3408_ (.A1(_0907_),
    .A2(\soc.cpu.AReg.data[8] ),
    .B1(_1012_),
    .B2(\soc.ram_data_out[8] ),
    .ZN(_1013_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3409_ (.A1(_1011_),
    .A2(_1013_),
    .ZN(_1014_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3410_ (.A1(_0853_),
    .A2(_1014_),
    .Z(_1015_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3411_ (.A1(_1010_),
    .A2(_1015_),
    .Z(_1016_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _3412_ (.A1(_1005_),
    .A2(_1008_),
    .A3(_1016_),
    .ZN(_1017_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3413_ (.A1(_0945_),
    .A2(_0981_),
    .A3(_1004_),
    .ZN(_1018_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _3414_ (.A1(_1000_),
    .A2(_1006_),
    .A3(_1007_),
    .ZN(_1019_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3415_ (.I(_1016_),
    .ZN(_1020_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3416_ (.A1(_1018_),
    .A2(_1019_),
    .B(_1020_),
    .ZN(_1021_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3417_ (.A1(_0875_),
    .A2(_1010_),
    .A3(_1015_),
    .ZN(_1022_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _3418_ (.A1(_0875_),
    .A2(_1017_),
    .A3(_1021_),
    .B(_1022_),
    .ZN(_1023_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3419_ (.A1(_0922_),
    .A2(_1023_),
    .ZN(_1024_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _3420_ (.A1(_0845_),
    .A2(_0926_),
    .B1(\soc.cpu.AReg.data[8] ),
    .B2(_0881_),
    .ZN(_1025_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3421_ (.A1(_0884_),
    .A2(_1024_),
    .B(_1025_),
    .ZN(\soc.cpu.PC.in[8] ));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3422_ (.A1(_1010_),
    .A2(_1015_),
    .ZN(_1026_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3423_ (.A1(_1005_),
    .A2(_1008_),
    .B(_1016_),
    .ZN(_1027_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3424_ (.A1(_0850_),
    .A2(\soc.cpu.ALU.x[9] ),
    .ZN(_1028_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3425_ (.A1(_0849_),
    .A2(_1028_),
    .ZN(_1029_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3426_ (.A1(_0907_),
    .A2(\soc.cpu.AReg.data[9] ),
    .B1(_1012_),
    .B2(\soc.ram_data_out[9] ),
    .ZN(_1030_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3427_ (.A1(_1011_),
    .A2(_1030_),
    .ZN(_1031_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3428_ (.A1(_0853_),
    .A2(_1031_),
    .Z(_1032_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3429_ (.A1(_1029_),
    .A2(_1032_),
    .Z(_1033_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3430_ (.I(_1033_),
    .ZN(_1034_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3431_ (.A1(_1026_),
    .A2(_1027_),
    .B(_1034_),
    .ZN(_1035_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _3432_ (.A1(_1026_),
    .A2(_1027_),
    .A3(_1034_),
    .Z(_1036_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3433_ (.A1(_0972_),
    .A2(_1029_),
    .A3(_1032_),
    .ZN(_1037_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _3434_ (.A1(_0972_),
    .A2(_1035_),
    .A3(_1036_),
    .B(_1037_),
    .ZN(_1038_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3435_ (.A1(_0990_),
    .A2(_1038_),
    .ZN(_1039_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _3436_ (.A1(_0845_),
    .A2(_1011_),
    .B1(\soc.cpu.AReg.data[9] ),
    .B2(_0880_),
    .ZN(_1040_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3437_ (.A1(_0884_),
    .A2(_1039_),
    .B(_1040_),
    .ZN(\soc.cpu.PC.in[9] ));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3438_ (.A1(_0904_),
    .A2(\soc.cpu.ALU.x[10] ),
    .ZN(_1041_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3439_ (.A1(_0923_),
    .A2(_1041_),
    .ZN(_1042_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3440_ (.A1(_0907_),
    .A2(\soc.cpu.AReg.data[10] ),
    .B1(_1012_),
    .B2(\soc.ram_data_out[10] ),
    .ZN(_1043_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3441_ (.A1(_1011_),
    .A2(_1043_),
    .ZN(_1044_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3442_ (.A1(_0926_),
    .A2(_1044_),
    .Z(_1045_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3443_ (.A1(_1042_),
    .A2(_1045_),
    .Z(_1046_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3444_ (.I(_1046_),
    .ZN(_1047_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3445_ (.A1(_1020_),
    .A2(_1034_),
    .ZN(_1048_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3446_ (.A1(_1005_),
    .A2(_1008_),
    .B(_1048_),
    .ZN(_1049_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3447_ (.A1(_1029_),
    .A2(_1032_),
    .ZN(_1050_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3448_ (.A1(_1029_),
    .A2(_1032_),
    .ZN(_1051_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3449_ (.A1(_1026_),
    .A2(_1050_),
    .B(_1051_),
    .ZN(_1052_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3450_ (.I(_1052_),
    .ZN(_1053_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _3451_ (.A1(_1047_),
    .A2(_1049_),
    .A3(_1053_),
    .Z(_1054_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3452_ (.A1(_1049_),
    .A2(_1053_),
    .B(_1047_),
    .ZN(_1055_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3453_ (.A1(_0972_),
    .A2(_1042_),
    .A3(_1045_),
    .ZN(_1056_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _3454_ (.A1(_0972_),
    .A2(_1054_),
    .A3(_1055_),
    .B(_1056_),
    .ZN(_1057_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3455_ (.A1(_0990_),
    .A2(_1057_),
    .ZN(_1058_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _3456_ (.A1(_0845_),
    .A2(_0923_),
    .B1(\soc.cpu.AReg.data[10] ),
    .B2(_0880_),
    .ZN(_1059_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3457_ (.A1(_0883_),
    .A2(_1058_),
    .B(_1059_),
    .ZN(\soc.cpu.PC.in[10] ));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _3458_ (.A1(_1042_),
    .A2(_1045_),
    .B(_1055_),
    .C(_0972_),
    .ZN(_1060_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3459_ (.A1(_0904_),
    .A2(\soc.cpu.ALU.x[11] ),
    .ZN(_1061_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3460_ (.A1(_0923_),
    .A2(_1061_),
    .ZN(_1062_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3461_ (.A1(_0907_),
    .A2(\soc.cpu.AReg.data[11] ),
    .B1(_1012_),
    .B2(\soc.ram_data_out[11] ),
    .ZN(_1063_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3462_ (.A1(_1011_),
    .A2(_1063_),
    .ZN(_1064_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3463_ (.A1(_0926_),
    .A2(_1064_),
    .Z(_1065_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3464_ (.A1(_1062_),
    .A2(_1065_),
    .ZN(_1066_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3465_ (.A1(_1062_),
    .A2(_1065_),
    .Z(_1067_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3466_ (.A1(_0954_),
    .A2(_1066_),
    .B(_1067_),
    .ZN(_1068_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _3467_ (.A1(_0922_),
    .A2(_1060_),
    .A3(_1068_),
    .Z(_1069_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _3468_ (.A1(_0846_),
    .A2(\soc.cpu.ALU.zx ),
    .B1(\soc.cpu.AReg.data[11] ),
    .B2(_0881_),
    .ZN(_1070_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3469_ (.A1(_0884_),
    .A2(_1069_),
    .B(_1070_),
    .ZN(\soc.cpu.PC.in[11] ));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3470_ (.A1(_0904_),
    .A2(\soc.cpu.ALU.x[12] ),
    .ZN(_1071_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3471_ (.A1(_0923_),
    .A2(_1071_),
    .ZN(_1072_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3472_ (.A1(_0907_),
    .A2(\soc.cpu.AReg.data[12] ),
    .B1(_1012_),
    .B2(\soc.ram_data_out[12] ),
    .ZN(_1073_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3473_ (.A1(_1011_),
    .A2(_1073_),
    .ZN(_1074_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3474_ (.A1(_0926_),
    .A2(_1074_),
    .Z(_1075_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3475_ (.A1(_1072_),
    .A2(_1075_),
    .ZN(_1076_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3476_ (.A1(_1067_),
    .A2(_1066_),
    .ZN(_1077_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3477_ (.A1(_1046_),
    .A2(_1048_),
    .A3(_1077_),
    .ZN(_1078_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3478_ (.I(_1078_),
    .ZN(_1079_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3479_ (.A1(_1005_),
    .A2(_1008_),
    .B(_1079_),
    .ZN(_1080_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3480_ (.A1(_1042_),
    .A2(_1045_),
    .ZN(_1081_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3481_ (.A1(_1046_),
    .A2(_1077_),
    .ZN(_1082_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _3482_ (.A1(_1081_),
    .A2(_1066_),
    .B1(_1082_),
    .B2(_1053_),
    .ZN(_1083_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3483_ (.A1(_1067_),
    .A2(_1083_),
    .ZN(_1084_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3484_ (.A1(_1072_),
    .A2(_1075_),
    .Z(_1085_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3485_ (.I(_1085_),
    .ZN(_1086_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _3486_ (.A1(_1080_),
    .A2(_1084_),
    .B(_1086_),
    .ZN(_1087_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3487_ (.A1(_1018_),
    .A2(_1019_),
    .B(_1078_),
    .ZN(_1088_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _3488_ (.A1(_1067_),
    .A2(_1083_),
    .Z(_1089_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _3489_ (.A1(_1088_),
    .A2(_1089_),
    .A3(_1085_),
    .B(_0954_),
    .ZN(_1090_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _3490_ (.A1(_0954_),
    .A2(_1076_),
    .B1(_1087_),
    .B2(_1090_),
    .ZN(_1091_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3491_ (.A1(_0990_),
    .A2(_1091_),
    .ZN(_1092_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _3492_ (.A1(_0845_),
    .A2(_0887_),
    .B1(\soc.cpu.AReg.data[12] ),
    .B2(_0880_),
    .ZN(_1093_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3493_ (.A1(_0883_),
    .A2(_1092_),
    .B(_1093_),
    .ZN(\soc.cpu.PC.in[12] ));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3494_ (.I(_1076_),
    .ZN(_1094_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3495_ (.A1(_0904_),
    .A2(\soc.cpu.ALU.x[13] ),
    .ZN(_1095_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3496_ (.A1(_0923_),
    .A2(_1095_),
    .ZN(_1096_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3497_ (.A1(_0907_),
    .A2(\soc.cpu.AReg.data[13] ),
    .B1(_1012_),
    .B2(\soc.ram_data_out[13] ),
    .ZN(_1097_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3498_ (.A1(_1011_),
    .A2(_1097_),
    .ZN(_1098_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3499_ (.A1(_0926_),
    .A2(_1098_),
    .Z(_1099_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3500_ (.A1(_1096_),
    .A2(_1099_),
    .Z(_1100_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _3501_ (.A1(_1094_),
    .A2(_1087_),
    .A3(_1100_),
    .ZN(_1101_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3502_ (.A1(_1088_),
    .A2(_1089_),
    .B(_1085_),
    .ZN(_1102_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3503_ (.I(_1100_),
    .ZN(_1103_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3504_ (.A1(_1076_),
    .A2(_1102_),
    .B(_1103_),
    .ZN(_1104_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3505_ (.A1(_1096_),
    .A2(_1099_),
    .Z(_1105_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3506_ (.A1(_0972_),
    .A2(_1105_),
    .ZN(_1106_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _3507_ (.A1(_0972_),
    .A2(_1101_),
    .A3(_1104_),
    .B(_1106_),
    .ZN(_1107_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _3508_ (.A1(_0990_),
    .A2(_1107_),
    .ZN(_1108_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _3509_ (.A1(_0845_),
    .A2(\soc.cpu.instruction[13] ),
    .B1(\soc.cpu.AReg.data[13] ),
    .B2(_0880_),
    .ZN(_1109_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3510_ (.A1(_0883_),
    .A2(_1108_),
    .B(_1109_),
    .ZN(\soc.cpu.PC.in[13] ));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3511_ (.A1(_0904_),
    .A2(\soc.cpu.ALU.x[14] ),
    .ZN(_1110_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3512_ (.A1(_0923_),
    .A2(_1110_),
    .ZN(_1111_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3513_ (.A1(_0907_),
    .A2(\soc.cpu.AReg.data[14] ),
    .B1(_1012_),
    .B2(\soc.ram_data_out[14] ),
    .ZN(_1112_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3514_ (.A1(_1011_),
    .A2(_1112_),
    .ZN(_1113_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3515_ (.A1(_0926_),
    .A2(_1113_),
    .Z(_1114_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3516_ (.A1(_1111_),
    .A2(_1114_),
    .Z(_1115_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _3517_ (.A1(_1105_),
    .A2(_1104_),
    .A3(_1115_),
    .ZN(_1116_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3518_ (.A1(_1096_),
    .A2(_1099_),
    .ZN(_1117_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3519_ (.A1(_1094_),
    .A2(_1087_),
    .B(_1100_),
    .ZN(_1118_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3520_ (.I(_1115_),
    .ZN(_1119_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3521_ (.A1(_1117_),
    .A2(_1118_),
    .B(_1119_),
    .ZN(_1120_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3522_ (.A1(_0972_),
    .A2(_1111_),
    .A3(_1114_),
    .ZN(_1121_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _3523_ (.A1(_0972_),
    .A2(_1116_),
    .A3(_1120_),
    .B(_1121_),
    .ZN(_1122_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3524_ (.A1(_0990_),
    .A2(_1122_),
    .ZN(_1123_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _3525_ (.A1(_0845_),
    .A2(\soc.cpu.instruction[14] ),
    .B1(\soc.cpu.AReg.data[14] ),
    .B2(_0880_),
    .ZN(_1124_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3526_ (.A1(_0883_),
    .A2(_1123_),
    .B(_1124_),
    .ZN(\soc.cpu.PC.in[14] ));
 gf180mcu_fd_sc_mcu7t5v0__inv_3 _3527_ (.I(\soc.video_generator_1.v_count[9] ),
    .ZN(_1125_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 _3528_ (.I(\soc.video_generator_1.v_count[6] ),
    .Z(_1126_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _3529_ (.I(\soc.video_generator_1.v_count[5] ),
    .Z(_1127_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _3530_ (.A1(\soc.video_generator_1.v_count[8] ),
    .A2(\soc.video_generator_1.v_count[7] ),
    .A3(_1126_),
    .A4(_1127_),
    .ZN(_1128_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3531_ (.A1(_1125_),
    .A2(_1128_),
    .ZN(_1129_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _3532_ (.I(\soc.video_generator_1.h_count[8] ),
    .ZN(_1130_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3533_ (.I(\soc.video_generator_1.h_count[6] ),
    .Z(_1131_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3534_ (.I(\soc.video_generator_1.h_count[7] ),
    .Z(_1132_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _3535_ (.A1(\soc.video_generator_1.h_count[5] ),
    .A2(_1131_),
    .B(_1132_),
    .ZN(_1133_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3536_ (.A1(_1130_),
    .A2(_1133_),
    .ZN(_1134_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3537_ (.A1(\soc.video_generator_1.h_count[9] ),
    .A2(_1134_),
    .ZN(_1135_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3538_ (.I(\soc.rom_encoder_0.initialized ),
    .ZN(_1136_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _3539_ (.A1(\soc.hack_wait_clocks[1] ),
    .A2(\soc.hack_wait_clocks[0] ),
    .A3(_1136_),
    .A4(_0741_),
    .ZN(_1137_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3540_ (.A1(\soc.ram_encoder_0.initialized ),
    .A2(\soc.spi_video_ram_1.initialized ),
    .A3(_1137_),
    .ZN(_1138_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _3541_ (.I(\soc.video_generator_1.v_count[0] ),
    .ZN(_1139_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _3542_ (.A1(_1125_),
    .A2(_1139_),
    .A3(_1128_),
    .ZN(_1140_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3543_ (.A1(\soc.boot_loading_offset[0] ),
    .A2(_1140_),
    .ZN(_1141_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 _3544_ (.I(\soc.video_generator_1.v_count[9] ),
    .Z(_1142_));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 _3545_ (.A1(\soc.video_generator_1.v_count[8] ),
    .A2(\soc.video_generator_1.v_count[7] ),
    .A3(\soc.video_generator_1.v_count[6] ),
    .A4(\soc.video_generator_1.v_count[5] ),
    .Z(_1143_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _3546_ (.A1(_1142_),
    .A2(\soc.video_generator_1.v_count[1] ),
    .A3(_1143_),
    .ZN(_1144_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3547_ (.A1(\soc.boot_loading_offset[1] ),
    .A2(_1144_),
    .ZN(_1145_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3548_ (.A1(\soc.boot_loading_offset[1] ),
    .A2(_1144_),
    .ZN(_1146_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _3549_ (.A1(_1141_),
    .A2(_1145_),
    .B(_1146_),
    .ZN(_1147_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3550_ (.A1(\soc.video_generator_1.v_count[2] ),
    .A2(\soc.video_generator_1.v_count[1] ),
    .ZN(_1148_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _3551_ (.A1(_1125_),
    .A2(_1128_),
    .A3(_1148_),
    .ZN(_1149_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _3552_ (.A1(_1142_),
    .A2(\soc.video_generator_1.v_count[2] ),
    .A3(\soc.video_generator_1.v_count[1] ),
    .A4(_1143_),
    .ZN(_1150_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _3553_ (.I(\soc.boot_loading_offset[2] ),
    .ZN(_1151_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _3554_ (.A1(_1149_),
    .A2(_1150_),
    .B(_1151_),
    .ZN(_1152_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _3555_ (.A1(_1151_),
    .A2(_1149_),
    .A3(_1150_),
    .ZN(_1153_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _3556_ (.A1(_1147_),
    .A2(_1152_),
    .B(_1153_),
    .C(\soc.boot_loading_offset[3] ),
    .ZN(_1154_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3557_ (.I(\soc.boot_loading_offset[3] ),
    .ZN(_1155_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _3558_ (.A1(_1149_),
    .A2(_1150_),
    .ZN(_1156_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3559_ (.A1(\soc.boot_loading_offset[2] ),
    .A2(_1156_),
    .ZN(_1157_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3560_ (.A1(\soc.boot_loading_offset[0] ),
    .A2(_1140_),
    .Z(_1158_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3561_ (.A1(\soc.boot_loading_offset[1] ),
    .A2(_1144_),
    .Z(_1159_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3562_ (.A1(\soc.boot_loading_offset[1] ),
    .A2(_1144_),
    .Z(_1160_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _3563_ (.A1(_1158_),
    .A2(_1159_),
    .B(_1153_),
    .C(_1160_),
    .ZN(_1161_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _3564_ (.I(\soc.video_generator_1.v_count[3] ),
    .ZN(_1162_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _3565_ (.A1(_1125_),
    .A2(_1162_),
    .A3(_1128_),
    .A4(_1148_),
    .ZN(_1163_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3566_ (.A1(\soc.video_generator_1.v_count[2] ),
    .A2(\soc.video_generator_1.v_count[1] ),
    .Z(_1164_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _3567_ (.A1(\soc.video_generator_1.v_count[3] ),
    .A2(_1164_),
    .B(_1143_),
    .C(_1142_),
    .ZN(_1165_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _3568_ (.A1(_1163_),
    .A2(_1165_),
    .Z(_1166_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 _3569_ (.I(\soc.video_generator_1.v_count[4] ),
    .Z(_1167_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _3570_ (.A1(\soc.video_generator_1.v_count[7] ),
    .A2(_1126_),
    .A3(_1127_),
    .ZN(_1168_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _3571_ (.A1(_1167_),
    .A2(_1168_),
    .ZN(_1169_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _3572_ (.A1(_1125_),
    .A2(_1139_),
    .A3(_1128_),
    .A4(_1164_),
    .ZN(_1170_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _3573_ (.A1(_1166_),
    .A2(_1169_),
    .A3(_1170_),
    .Z(_1171_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _3574_ (.A1(_1155_),
    .A2(_1157_),
    .A3(_1161_),
    .B(_1171_),
    .ZN(_1172_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3575_ (.A1(_1166_),
    .A2(_1169_),
    .ZN(_1173_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _3576_ (.A1(\soc.boot_loading_offset[2] ),
    .A2(_1156_),
    .A3(_1147_),
    .Z(_1174_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _3577_ (.A1(_1173_),
    .A2(_1156_),
    .B1(_1171_),
    .B2(_1174_),
    .ZN(_1175_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _3578_ (.A1(_1154_),
    .A2(_1172_),
    .B(_1166_),
    .C(_1175_),
    .ZN(_1176_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3579_ (.A1(_1163_),
    .A2(_1165_),
    .ZN(_1177_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3580_ (.A1(\soc.boot_loading_offset[3] ),
    .A2(_1177_),
    .ZN(_1178_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3581_ (.A1(\soc.boot_loading_offset[3] ),
    .A2(_1177_),
    .ZN(_1179_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _3582_ (.A1(_1157_),
    .A2(_1161_),
    .A3(_1178_),
    .B(_1179_),
    .ZN(_1180_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3583_ (.A1(\soc.video_generator_1.v_count[4] ),
    .A2(_1129_),
    .ZN(_1181_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3584_ (.I0(\soc.video_generator_1.v_count[4] ),
    .I1(_1181_),
    .S(_1163_),
    .Z(_1182_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3585_ (.A1(\soc.boot_loading_offset[4] ),
    .A2(_1182_),
    .ZN(_1183_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3586_ (.A1(_1180_),
    .A2(_1183_),
    .Z(_1184_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3587_ (.A1(_1180_),
    .A2(_1183_),
    .B(_1171_),
    .ZN(_1185_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _3588_ (.A1(_1184_),
    .A2(_1185_),
    .B(_1182_),
    .ZN(_1186_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3589_ (.A1(_1130_),
    .A2(\soc.video_generator_1.h_count[9] ),
    .A3(_1133_),
    .ZN(_1187_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _3590_ (.A1(_1130_),
    .A2(_1133_),
    .B(_1187_),
    .ZN(_1188_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _3591_ (.A1(\soc.video_generator_1.h_count[8] ),
    .A2(\soc.video_generator_1.h_count[9] ),
    .ZN(_1189_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3592_ (.I(\soc.video_generator_1.h_count[5] ),
    .Z(_1190_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _3593_ (.A1(_1190_),
    .A2(_1132_),
    .A3(_1131_),
    .ZN(_1191_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3594_ (.A1(_1189_),
    .A2(_1191_),
    .ZN(_1192_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3595_ (.A1(_1133_),
    .A2(_1192_),
    .ZN(_1193_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3596_ (.A1(\soc.video_generator_1.h_count[5] ),
    .A2(_1131_),
    .Z(_1194_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _3597_ (.A1(_1135_),
    .A2(_1194_),
    .Z(_1195_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _3598_ (.A1(_1133_),
    .A2(_1189_),
    .ZN(_1196_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3599_ (.A1(\soc.video_generator_1.h_count[3] ),
    .A2(\soc.video_generator_1.h_count[4] ),
    .A3(_1196_),
    .ZN(_1197_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _3600_ (.A1(\soc.video_generator_1.h_count[5] ),
    .A2(_1197_),
    .Z(_1198_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3601_ (.A1(_1195_),
    .A2(_1198_),
    .Z(_1199_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3602_ (.A1(_1193_),
    .A2(_1199_),
    .ZN(_1200_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3603_ (.A1(_1188_),
    .A2(_1200_),
    .Z(_1201_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _3604_ (.A1(_1176_),
    .A2(_1186_),
    .A3(_1201_),
    .ZN(_1202_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3605_ (.A1(_1193_),
    .A2(_1199_),
    .Z(_1203_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3606_ (.A1(_1154_),
    .A2(_1172_),
    .B(_1166_),
    .ZN(_1204_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3607_ (.A1(_1175_),
    .A2(_1204_),
    .ZN(_1205_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3608_ (.A1(_1203_),
    .A2(_1205_),
    .ZN(_1206_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _3609_ (.A1(\soc.video_generator_1.h_count[3] ),
    .A2(\soc.video_generator_1.h_count[4] ),
    .Z(_1207_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _3610_ (.A1(_1196_),
    .A2(_1197_),
    .A3(_1207_),
    .Z(_1208_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3611_ (.I(\soc.boot_loading_offset[0] ),
    .ZN(_1209_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _3612_ (.A1(_1163_),
    .A2(_1165_),
    .A3(_1169_),
    .A4(_1170_),
    .ZN(_1210_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _3613_ (.A1(_1142_),
    .A2(_1143_),
    .ZN(_1211_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _3614_ (.A1(_1209_),
    .A2(_1210_),
    .B(_1211_),
    .C(_1139_),
    .ZN(_1212_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _3615_ (.A1(_1166_),
    .A2(_1169_),
    .A3(_1158_),
    .ZN(_1213_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3616_ (.A1(_1208_),
    .A2(_1212_),
    .A3(_1213_),
    .ZN(_1214_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3617_ (.A1(\soc.video_generator_1.h_count[3] ),
    .A2(_1196_),
    .ZN(_1215_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3618_ (.I(\soc.display_clks_before_active[0] ),
    .Z(_1216_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _3619_ (.A1(_1216_),
    .A2(_1196_),
    .ZN(_1217_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3620_ (.A1(\soc.video_generator_1.h_count[1] ),
    .A2(_1196_),
    .ZN(_1218_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3621_ (.A1(\soc.video_generator_1.h_count[2] ),
    .A2(_1196_),
    .ZN(_1219_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _3622_ (.A1(_1217_),
    .A2(_1218_),
    .A3(_1219_),
    .ZN(_1220_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3623_ (.A1(_1215_),
    .A2(_1220_),
    .ZN(_1221_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _3624_ (.A1(_1212_),
    .A2(_1213_),
    .B(_1208_),
    .ZN(_1222_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _3625_ (.A1(_1214_),
    .A2(_1221_),
    .B(_1222_),
    .ZN(_1223_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3626_ (.A1(_1158_),
    .A2(_1159_),
    .Z(_1224_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3627_ (.A1(_1144_),
    .A2(_1173_),
    .B1(_1171_),
    .B2(_1224_),
    .ZN(_1225_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3628_ (.A1(_1190_),
    .A2(_1135_),
    .B(_1197_),
    .ZN(_1226_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3629_ (.A1(_1198_),
    .A2(_1226_),
    .ZN(_1227_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3630_ (.A1(_1225_),
    .A2(_1227_),
    .ZN(_1228_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3631_ (.A1(_1225_),
    .A2(_1227_),
    .ZN(_1229_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _3632_ (.A1(_1223_),
    .A2(_1228_),
    .B(_1229_),
    .ZN(_1230_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3633_ (.A1(_1195_),
    .A2(_1198_),
    .ZN(_1231_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3634_ (.A1(_1175_),
    .A2(_1231_),
    .Z(_1232_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3635_ (.A1(_1175_),
    .A2(_1231_),
    .ZN(_1233_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _3636_ (.A1(_1203_),
    .A2(_1205_),
    .B1(_1230_),
    .B2(_1232_),
    .C(_1233_),
    .ZN(_1234_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3637_ (.A1(_1206_),
    .A2(_1234_),
    .ZN(_1235_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3638_ (.A1(_1202_),
    .A2(_1235_),
    .ZN(_1236_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3639_ (.A1(_1230_),
    .A2(_1232_),
    .B(_1233_),
    .ZN(_1237_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _3640_ (.A1(_1203_),
    .A2(_1205_),
    .A3(_1237_),
    .Z(_1238_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _3641_ (.A1(_1223_),
    .A2(_1228_),
    .ZN(_1239_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _3642_ (.A1(_1208_),
    .A2(_1212_),
    .A3(_1213_),
    .Z(_1240_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _3643_ (.A1(_1222_),
    .A2(_1240_),
    .ZN(_1241_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3644_ (.A1(_1127_),
    .A2(_1211_),
    .ZN(_1242_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _3645_ (.A1(_1167_),
    .A2(_1163_),
    .Z(_1243_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3646_ (.A1(_1242_),
    .A2(_1243_),
    .Z(_1244_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3647_ (.A1(_1171_),
    .A2(_1180_),
    .A3(_1183_),
    .ZN(_1245_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3648_ (.A1(_1244_),
    .A2(_1245_),
    .ZN(_1246_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _3649_ (.A1(_1176_),
    .A2(_1186_),
    .B(_1246_),
    .ZN(_1247_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _3650_ (.A1(_1176_),
    .A2(_1186_),
    .A3(_1246_),
    .Z(_1248_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3651_ (.A1(\soc.video_generator_1.h_count[9] ),
    .A2(_1134_),
    .ZN(_1249_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3652_ (.A1(_1188_),
    .A2(_1200_),
    .ZN(_1250_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3653_ (.A1(_1249_),
    .A2(_1250_),
    .ZN(_1251_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3654_ (.A1(_1247_),
    .A2(_1248_),
    .B(_1251_),
    .ZN(_1252_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3655_ (.A1(_1176_),
    .A2(_1186_),
    .Z(_1253_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _3656_ (.A1(_1202_),
    .A2(_1206_),
    .A3(_1234_),
    .B1(_1201_),
    .B2(_1253_),
    .ZN(_1254_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _3657_ (.A1(_1247_),
    .A2(_1248_),
    .A3(_1251_),
    .ZN(_1255_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3658_ (.A1(_1252_),
    .A2(_1254_),
    .B(_1255_),
    .ZN(_1256_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3659_ (.A1(_1142_),
    .A2(_1126_),
    .ZN(_1257_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3660_ (.A1(_1127_),
    .A2(_1211_),
    .A3(_1243_),
    .ZN(_1258_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3661_ (.I0(_1126_),
    .I1(_1257_),
    .S(_1258_),
    .Z(_1259_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _3662_ (.A1(_1247_),
    .A2(_1256_),
    .A3(_1259_),
    .Z(_1260_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3663_ (.I(_1260_),
    .Z(_1261_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _3664_ (.A1(\soc.video_generator_1.h_count[1] ),
    .A2(\soc.video_generator_1.h_count[2] ),
    .A3(_1215_),
    .ZN(_1262_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _3665_ (.A1(_1241_),
    .A2(_1261_),
    .A3(_1262_),
    .ZN(_1263_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3666_ (.A1(_1239_),
    .A2(_1263_),
    .ZN(_1264_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3667_ (.A1(_1215_),
    .A2(_1220_),
    .ZN(_1265_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3668_ (.A1(\soc.video_generator_1.h_count[2] ),
    .A2(_1217_),
    .ZN(_1266_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3669_ (.A1(_1218_),
    .A2(_1266_),
    .B(_1261_),
    .ZN(_1267_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3670_ (.A1(\soc.video_generator_1.h_count[1] ),
    .A2(_1216_),
    .ZN(_1268_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3671_ (.A1(_1268_),
    .A2(_1219_),
    .B(_1220_),
    .ZN(_1269_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3672_ (.A1(_1217_),
    .A2(_1269_),
    .Z(_1270_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3673_ (.A1(_1261_),
    .A2(_1270_),
    .B(_1265_),
    .ZN(_1271_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3674_ (.A1(_1241_),
    .A2(_1221_),
    .Z(_1272_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3675_ (.A1(_1265_),
    .A2(_1267_),
    .B(_1271_),
    .C(_1272_),
    .ZN(_1273_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3676_ (.A1(_1261_),
    .A2(_1262_),
    .ZN(_1274_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3677_ (.A1(_1241_),
    .A2(_1274_),
    .ZN(_1275_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3678_ (.A1(_1230_),
    .A2(_1232_),
    .ZN(_1276_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _3679_ (.A1(_1264_),
    .A2(_1273_),
    .B1(_1275_),
    .B2(_1239_),
    .C(_1276_),
    .ZN(_1277_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3680_ (.A1(_1217_),
    .A2(_1218_),
    .ZN(_1278_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3681_ (.I(_1272_),
    .ZN(_1279_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _3682_ (.I(_1239_),
    .ZN(_1280_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3683_ (.A1(\soc.video_generator_1.h_count[1] ),
    .A2(_1216_),
    .Z(_1281_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3684_ (.A1(_1279_),
    .A2(_1280_),
    .A3(_1281_),
    .ZN(_1282_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3685_ (.A1(_1272_),
    .A2(_1239_),
    .B(_1270_),
    .ZN(_1283_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3686_ (.A1(_1272_),
    .A2(_1239_),
    .A3(_1266_),
    .ZN(_1284_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _3687_ (.A1(_1278_),
    .A2(_1282_),
    .A3(_1283_),
    .A4(_1284_),
    .ZN(_1285_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _3688_ (.A1(_1215_),
    .A2(_1220_),
    .Z(_1286_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3689_ (.A1(_1196_),
    .A2(_1281_),
    .ZN(_1287_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3690_ (.A1(_1278_),
    .A2(_1287_),
    .ZN(_1288_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3691_ (.A1(_1241_),
    .A2(_1288_),
    .ZN(_1289_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3692_ (.A1(_1286_),
    .A2(_1280_),
    .ZN(_1290_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3693_ (.A1(_1288_),
    .A2(_1290_),
    .B(_1269_),
    .ZN(_1291_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3694_ (.A1(_1286_),
    .A2(_1289_),
    .B(_1291_),
    .ZN(_1292_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3695_ (.A1(_1217_),
    .A2(_1292_),
    .B(_1276_),
    .ZN(_1293_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _3696_ (.A1(_1265_),
    .A2(_1285_),
    .B(_1293_),
    .C(_1261_),
    .ZN(_1294_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3697_ (.A1(_1277_),
    .A2(_1294_),
    .ZN(_1295_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3698_ (.A1(\soc.video_generator_1.h_count[3] ),
    .A2(\soc.video_generator_1.h_count[2] ),
    .ZN(_1296_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3699_ (.A1(\soc.video_generator_1.h_count[1] ),
    .A2(_1216_),
    .B(_1218_),
    .ZN(_1297_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3700_ (.A1(_1216_),
    .A2(_1218_),
    .B(_1219_),
    .ZN(_1298_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3701_ (.A1(_1297_),
    .A2(_1298_),
    .ZN(_1299_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3702_ (.A1(_1278_),
    .A2(_1296_),
    .B1(_1299_),
    .B2(_1286_),
    .ZN(_1300_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3703_ (.A1(\soc.video_generator_1.h_count[3] ),
    .A2(_1196_),
    .B(_1269_),
    .ZN(_1301_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3704_ (.A1(_1280_),
    .A2(_1301_),
    .A3(_1288_),
    .ZN(_1302_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _3705_ (.A1(_1280_),
    .A2(_1300_),
    .B1(_1290_),
    .B2(_1217_),
    .C(_1302_),
    .ZN(_1303_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3706_ (.A1(_1286_),
    .A2(_1261_),
    .B(_1303_),
    .ZN(_1304_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3707_ (.A1(_1271_),
    .A2(_1304_),
    .ZN(_1305_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _3708_ (.A1(_1260_),
    .A2(_1301_),
    .A3(_1287_),
    .B(_1265_),
    .ZN(_1306_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _3709_ (.A1(_1216_),
    .A2(\soc.video_generator_1.h_count[2] ),
    .A3(_1218_),
    .Z(_1307_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3710_ (.A1(_1261_),
    .A2(_1307_),
    .B(_1286_),
    .ZN(_1308_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3711_ (.A1(_1306_),
    .A2(_1308_),
    .B(_1279_),
    .ZN(_1309_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _3712_ (.A1(_1279_),
    .A2(_1305_),
    .B(_1309_),
    .C(_1276_),
    .ZN(_1310_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3713_ (.I(_1276_),
    .ZN(_1311_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3714_ (.A1(_1286_),
    .A2(_1269_),
    .B(_1301_),
    .ZN(_1312_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3715_ (.A1(_1261_),
    .A2(_1312_),
    .B(_1239_),
    .ZN(_1313_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3716_ (.A1(_1272_),
    .A2(_1313_),
    .B(_1263_),
    .ZN(_1314_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _3717_ (.A1(_1280_),
    .A2(_1309_),
    .B(_1311_),
    .C(_1314_),
    .ZN(_1315_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _3718_ (.A1(_1310_),
    .A2(_1238_),
    .A3(_1315_),
    .ZN(_1316_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3719_ (.A1(_1238_),
    .A2(_1295_),
    .B(_1316_),
    .ZN(_1317_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _3720_ (.A1(_1236_),
    .A2(_1317_),
    .Z(_1318_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3721_ (.A1(_1261_),
    .A2(_1307_),
    .ZN(_1319_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3722_ (.A1(_1261_),
    .A2(_1266_),
    .B(_1279_),
    .C(_1286_),
    .ZN(_1320_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3723_ (.A1(_1306_),
    .A2(_1319_),
    .B(_1320_),
    .ZN(_1321_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3724_ (.A1(_1309_),
    .A2(_1321_),
    .B(_1239_),
    .ZN(_1322_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3725_ (.A1(_1311_),
    .A2(_1264_),
    .ZN(_1323_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3726_ (.A1(_1238_),
    .A2(_1322_),
    .A3(_1323_),
    .ZN(_1324_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3727_ (.A1(_1236_),
    .A2(_1324_),
    .ZN(_1325_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3728_ (.A1(_1193_),
    .A2(_1195_),
    .ZN(_1326_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3729_ (.A1(\soc.video_generator_1.h_count[3] ),
    .A2(_1196_),
    .A3(_1220_),
    .ZN(_1327_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3730_ (.I(_1132_),
    .ZN(_1328_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3731_ (.A1(\soc.video_generator_1.h_count[4] ),
    .A2(_1328_),
    .ZN(_1329_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _3732_ (.A1(_1190_),
    .A2(_1131_),
    .A3(_1327_),
    .A4(_1329_),
    .ZN(_1330_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3733_ (.A1(\soc.video_generator_1.v_count[3] ),
    .A2(_1129_),
    .ZN(_1331_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _3734_ (.A1(_1331_),
    .A2(_1150_),
    .A3(_1181_),
    .ZN(_1332_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3735_ (.I(_1126_),
    .ZN(_1333_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3736_ (.A1(_1142_),
    .A2(\soc.video_generator_1.v_count[7] ),
    .B(_1249_),
    .C(_1188_),
    .ZN(_1334_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _3737_ (.A1(_1333_),
    .A2(_1242_),
    .A3(_1208_),
    .A4(_1334_),
    .ZN(_1335_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3738_ (.A1(_1162_),
    .A2(\soc.video_generator_1.v_count[2] ),
    .ZN(_1336_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3739_ (.A1(_1167_),
    .A2(_1336_),
    .ZN(_1337_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _3740_ (.A1(\soc.video_generator_1.v_count[1] ),
    .A2(_1168_),
    .A3(_1129_),
    .A4(_1337_),
    .ZN(_1338_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3741_ (.A1(_1140_),
    .A2(_1338_),
    .B(_1199_),
    .ZN(_1339_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3742_ (.A1(_1243_),
    .A2(_1335_),
    .A3(_1339_),
    .ZN(_1340_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _3743_ (.A1(_1326_),
    .A2(_1330_),
    .B(_1332_),
    .C(_1340_),
    .ZN(_1341_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3744_ (.A1(_1247_),
    .A2(_1248_),
    .ZN(_1342_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _3745_ (.A1(_1342_),
    .A2(_1251_),
    .A3(_1254_),
    .Z(_1343_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _3746_ (.A1(_1318_),
    .A2(_1325_),
    .A3(_1341_),
    .A4(_1343_),
    .ZN(_1344_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3747_ (.A1(_1196_),
    .A2(_1249_),
    .ZN(_1345_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _3748_ (.A1(_1326_),
    .A2(_1188_),
    .Z(_1346_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3749_ (.I0(\soc.spi_video_ram_1.read_value[2] ),
    .I1(\soc.spi_video_ram_1.read_value[3] ),
    .S(_1217_),
    .Z(_1347_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _3750_ (.A1(_1345_),
    .A2(_1346_),
    .B1(_1218_),
    .B2(_1347_),
    .C(_1138_),
    .ZN(_1348_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3751_ (.I(\soc.spi_video_ram_1.read_value[1] ),
    .ZN(_1349_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3752_ (.A1(\soc.spi_video_ram_1.read_value[0] ),
    .A2(_1217_),
    .ZN(_1350_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _3753_ (.A1(_1349_),
    .A2(_1217_),
    .B(_1218_),
    .C(_1350_),
    .ZN(_1351_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3754_ (.A1(_1142_),
    .A2(\soc.video_generator_1.v_count[8] ),
    .ZN(_1352_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _3755_ (.A1(_1142_),
    .A2(\soc.video_generator_1.v_count[7] ),
    .ZN(_1353_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _3756_ (.A1(_1126_),
    .A2(_1127_),
    .A3(_1167_),
    .A4(_1211_),
    .ZN(_1354_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3757_ (.A1(_1353_),
    .A2(_1354_),
    .ZN(_1355_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3758_ (.A1(_1352_),
    .A2(_1355_),
    .Z(_1356_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _3759_ (.A1(_1189_),
    .A2(_1195_),
    .B(_1351_),
    .C(_1356_),
    .ZN(_1357_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3760_ (.A1(_1138_),
    .A2(_1344_),
    .B1(_1348_),
    .B2(_1357_),
    .ZN(_1358_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _3761_ (.A1(_1129_),
    .A2(_1135_),
    .A3(_1358_),
    .ZN(net76));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _3762_ (.I(\soc.ram_encoder_0.sram_sio_oe ),
    .ZN(net49));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _3763_ (.I(\soc.rom_encoder_0.sram_sio_oe ),
    .ZN(net53));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _3764_ (.I(\soc.spi_video_ram_1.sram_sio_oe ),
    .ZN(net57));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3765_ (.A1(\soc.video_generator_1.h_count[4] ),
    .A2(_1190_),
    .A3(_1131_),
    .ZN(_1359_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _3766_ (.A1(\soc.video_generator_1.h_count[4] ),
    .A2(_1190_),
    .A3(_1131_),
    .Z(_1360_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _3767_ (.A1(_1328_),
    .A2(_1189_),
    .A3(_1359_),
    .A4(_1360_),
    .ZN(net75));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3768_ (.A1(\soc.video_generator_1.v_count[8] ),
    .A2(\soc.video_generator_1.v_count[1] ),
    .Z(_1361_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _3769_ (.A1(_1125_),
    .A2(_1169_),
    .A3(_1336_),
    .A4(_1361_),
    .ZN(net74));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3770_ (.A1(_0752_),
    .A2(_0808_),
    .Z(_1362_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _3771_ (.A1(_0758_),
    .A2(_0759_),
    .A3(_0752_),
    .ZN(_1363_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3772_ (.A1(_0749_),
    .A2(_1363_),
    .Z(_1364_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3773_ (.A1(_0760_),
    .A2(_0830_),
    .ZN(_1365_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3774_ (.A1(_0811_),
    .A2(_0825_),
    .B1(_0827_),
    .B2(_0815_),
    .ZN(_1366_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3775_ (.A1(_1365_),
    .A2(_1366_),
    .ZN(_1367_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _3776_ (.A1(_0808_),
    .A2(_0822_),
    .B(_1364_),
    .C(_1367_),
    .ZN(_1368_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _3777_ (.A1(_0776_),
    .A2(\soc.spi_video_ram_1.output_buffer[1] ),
    .A3(_0811_),
    .Z(_1369_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3778_ (.A1(_0808_),
    .A2(_0838_),
    .B(_0760_),
    .ZN(_1370_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3779_ (.A1(_0836_),
    .A2(_1370_),
    .B(_1364_),
    .ZN(_1371_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _3780_ (.A1(_0815_),
    .A2(_0839_),
    .B(_1369_),
    .C(_1371_),
    .ZN(_1372_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3781_ (.A1(_0808_),
    .A2(_0814_),
    .B1(_0816_),
    .B2(_0760_),
    .ZN(_1373_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3782_ (.A1(_0771_),
    .A2(_1373_),
    .ZN(_1374_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _3783_ (.A1(_0809_),
    .A2(_0811_),
    .B1(_0812_),
    .B2(_0815_),
    .C(_1374_),
    .ZN(_1375_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3784_ (.A1(_1364_),
    .A2(_1362_),
    .ZN(_1376_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _3785_ (.A1(_1362_),
    .A2(_1368_),
    .A3(_1372_),
    .B1(_1375_),
    .B2(_1376_),
    .ZN(_1377_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3786_ (.A1(_0807_),
    .A2(_1377_),
    .Z(_1378_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3787_ (.I(_1378_),
    .Z(net71));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3788_ (.A1(_0759_),
    .A2(_0763_),
    .Z(_1379_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3789_ (.A1(_0775_),
    .A2(_0790_),
    .ZN(_1380_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3790_ (.A1(_0775_),
    .A2(_0787_),
    .B(_1379_),
    .C(_1380_),
    .ZN(_1381_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3791_ (.A1(_0763_),
    .A2(_0753_),
    .ZN(_1382_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _3792_ (.A1(\soc.spi_video_ram_1.buffer_index[4] ),
    .A2(_1382_),
    .Z(_1383_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _3793_ (.A1(_0779_),
    .A2(_0784_),
    .B1(_0785_),
    .B2(_0765_),
    .C(_1379_),
    .ZN(_1384_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3794_ (.A1(_0759_),
    .A2(_0764_),
    .B(_0752_),
    .ZN(_1385_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3795_ (.A1(_1382_),
    .A2(_1385_),
    .Z(_1386_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3796_ (.A1(_1384_),
    .A2(_1386_),
    .ZN(_1387_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3797_ (.A1(_1381_),
    .A2(_1383_),
    .A3(_1387_),
    .ZN(_1388_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3798_ (.I0(\soc.spi_video_ram_1.output_buffer[19] ),
    .I1(\soc.spi_video_ram_1.output_buffer[16] ),
    .I2(\soc.spi_video_ram_1.output_buffer[17] ),
    .I3(\soc.spi_video_ram_1.output_buffer[18] ),
    .S0(_0757_),
    .S1(_0758_),
    .Z(_1389_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3799_ (.I(_1389_),
    .ZN(_1390_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3800_ (.A1(_0758_),
    .A2(\soc.spi_video_ram_1.output_buffer[1] ),
    .B(_0775_),
    .ZN(_1391_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3801_ (.A1(_0761_),
    .A2(_0766_),
    .B(_1383_),
    .ZN(_1392_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _3802_ (.A1(_1383_),
    .A2(_1390_),
    .B1(_1391_),
    .B2(_1392_),
    .ZN(_1393_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3803_ (.I0(_0794_),
    .I1(_0796_),
    .S(_0765_),
    .Z(_1394_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3804_ (.A1(_0765_),
    .A2(_0777_),
    .ZN(_1395_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3805_ (.A1(_0775_),
    .A2(_0773_),
    .ZN(_1396_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3806_ (.A1(_1383_),
    .A2(_1395_),
    .A3(_1396_),
    .ZN(_1397_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3807_ (.A1(_1383_),
    .A2(_1394_),
    .B(_1397_),
    .C(_1379_),
    .ZN(_1398_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3808_ (.A1(_1379_),
    .A2(_1393_),
    .B(_1398_),
    .C(_1386_),
    .ZN(_1399_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3809_ (.A1(\soc.spi_video_ram_1.buffer_index[4] ),
    .A2(_1382_),
    .B(\soc.spi_video_ram_1.buffer_index[5] ),
    .ZN(_1400_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3810_ (.A1(_0764_),
    .A2(_0770_),
    .B(_1400_),
    .ZN(_1401_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _3811_ (.A1(_1388_),
    .A2(_1399_),
    .B(_1401_),
    .C(_0720_),
    .ZN(net72));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _3812_ (.A1(_0720_),
    .A2(_0843_),
    .Z(_1402_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3813_ (.I(_1402_),
    .Z(net73));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3814_ (.I(\soc.rom_encoder_0.toggled_sram_sck ),
    .Z(_1403_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3815_ (.I(_1403_),
    .ZN(_1404_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3816_ (.A1(net62),
    .A2(_1404_),
    .ZN(net63));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3817_ (.I(\soc.ram_encoder_0.toggled_sram_sck ),
    .ZN(_1405_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3818_ (.A1(net81),
    .A2(_1405_),
    .ZN(net82));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _3819_ (.I(\soc.rom_encoder_0.current_state[0] ),
    .Z(_1406_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_3 _3820_ (.I(\soc.rom_encoder_0.current_state[2] ),
    .ZN(_1407_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _3821_ (.I(\soc.rom_encoder_0.current_state[1] ),
    .ZN(_1408_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3822_ (.A1(_1407_),
    .A2(_1408_),
    .ZN(_1409_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3823_ (.A1(_1406_),
    .A2(_1409_),
    .ZN(_1410_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3824_ (.I(\soc.rom_encoder_0.request_write ),
    .ZN(_1411_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _3825_ (.A1(\soc.rom_encoder_0.current_state[2] ),
    .A2(_1408_),
    .ZN(_1412_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3826_ (.A1(_1406_),
    .A2(_1412_),
    .ZN(_1413_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3827_ (.I(\soc.rom_encoder_0.output_bits_left[4] ),
    .ZN(_1414_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3828_ (.I(\soc.rom_encoder_0.output_bits_left[3] ),
    .ZN(_1415_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3829_ (.A1(\soc.rom_encoder_0.output_bits_left[2] ),
    .A2(_1414_),
    .A3(_1415_),
    .ZN(_1416_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _3830_ (.I(_1416_),
    .Z(_1417_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3831_ (.A1(_1413_),
    .A2(_1417_),
    .ZN(_1418_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _3832_ (.I(_1406_),
    .ZN(_1419_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3833_ (.A1(\soc.rom_encoder_0.current_state[1] ),
    .A2(_1419_),
    .ZN(_1420_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3834_ (.A1(\soc.rom_encoder_0.current_state[2] ),
    .A2(_1420_),
    .ZN(_1421_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3835_ (.A1(_1408_),
    .A2(_1419_),
    .ZN(_1422_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3836_ (.A1(_1416_),
    .A2(_1421_),
    .B(_1422_),
    .C(_1403_),
    .ZN(_1423_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _3837_ (.A1(_1411_),
    .A2(_1418_),
    .B(_1423_),
    .ZN(_1424_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _3838_ (.A1(\soc.rom_encoder_0.initializing_step[4] ),
    .A2(\soc.rom_encoder_0.initializing_step[3] ),
    .A3(\soc.rom_encoder_0.initializing_step[2] ),
    .A4(\soc.rom_encoder_0.initializing_step[1] ),
    .Z(_1425_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3839_ (.I(\soc.rom_encoder_0.current_state[2] ),
    .Z(_1426_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3840_ (.A1(_1426_),
    .A2(\soc.rom_encoder_0.current_state[1] ),
    .ZN(_1427_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3841_ (.A1(_1406_),
    .A2(_1427_),
    .ZN(_1428_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3842_ (.A1(_1425_),
    .A2(_1428_),
    .ZN(_1429_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3843_ (.A1(_1424_),
    .A2(_1429_),
    .ZN(_1430_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _3844_ (.I(_1430_),
    .ZN(_1431_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3845_ (.A1(_1410_),
    .A2(_1431_),
    .ZN(_1432_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3846_ (.A1(\soc.rom_encoder_0.output_bits_left[2] ),
    .A2(_1415_),
    .ZN(_1433_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _3847_ (.A1(\soc.rom_encoder_0.output_bits_left[4] ),
    .A2(_1433_),
    .ZN(_1434_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3848_ (.A1(_1426_),
    .A2(_1419_),
    .ZN(_1435_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _3849_ (.A1(_1412_),
    .A2(_1434_),
    .B(_1435_),
    .ZN(_1436_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3850_ (.A1(_1427_),
    .A2(_1422_),
    .ZN(_1437_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3851_ (.I(\soc.rom_encoder_0.initializing_step[0] ),
    .Z(_1438_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _3852_ (.A1(\soc.rom_encoder_0.initializing_step[4] ),
    .A2(\soc.rom_encoder_0.initializing_step[3] ),
    .A3(\soc.rom_encoder_0.initializing_step[2] ),
    .A4(\soc.rom_encoder_0.initializing_step[1] ),
    .ZN(_1439_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3853_ (.A1(_1438_),
    .A2(_1439_),
    .ZN(_1440_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3854_ (.A1(_1437_),
    .A2(_1440_),
    .Z(_1441_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _3855_ (.A1(_1417_),
    .A2(_1437_),
    .ZN(_1442_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3856_ (.A1(\soc.rom_encoder_0.output_buffer[17] ),
    .A2(_1417_),
    .B1(_1442_),
    .B2(\soc.rom_encoder_0.request_data_out[13] ),
    .ZN(_1443_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3857_ (.A1(_1413_),
    .A2(_1443_),
    .ZN(_1444_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _3858_ (.A1(\soc.rom_encoder_0.output_buffer[17] ),
    .A2(_1436_),
    .B(_1441_),
    .C(_1444_),
    .ZN(_1445_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3859_ (.A1(net65),
    .A2(_1432_),
    .ZN(_1446_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3860_ (.A1(_1432_),
    .A2(_1445_),
    .B(_1446_),
    .C(_0676_),
    .ZN(_0010_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3861_ (.A1(\soc.rom_encoder_0.output_buffer[18] ),
    .A2(_1417_),
    .B1(_1442_),
    .B2(\soc.rom_encoder_0.request_data_out[14] ),
    .ZN(_1447_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3862_ (.A1(_1413_),
    .A2(_1447_),
    .ZN(_1448_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _3863_ (.A1(\soc.rom_encoder_0.output_buffer[18] ),
    .A2(_1436_),
    .B(_1448_),
    .C(_1441_),
    .ZN(_1449_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3864_ (.A1(net66),
    .A2(_1432_),
    .ZN(_1450_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3865_ (.A1(_1432_),
    .A2(_1449_),
    .B(_1450_),
    .C(_0676_),
    .ZN(_0011_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3866_ (.A1(\soc.rom_encoder_0.output_buffer[19] ),
    .A2(_1417_),
    .B1(_1442_),
    .B2(\soc.rom_encoder_0.request_data_out[15] ),
    .ZN(_1451_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3867_ (.A1(_1413_),
    .A2(_1451_),
    .ZN(_1452_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _3868_ (.A1(\soc.rom_encoder_0.output_buffer[19] ),
    .A2(_1436_),
    .B(_1452_),
    .C(_1441_),
    .ZN(_1453_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3869_ (.A1(net67),
    .A2(_1432_),
    .ZN(_1454_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3870_ (.A1(_1432_),
    .A2(_1453_),
    .B(_1454_),
    .C(_0676_),
    .ZN(_0012_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3871_ (.A1(_1190_),
    .A2(_1296_),
    .ZN(_1455_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3872_ (.A1(\soc.video_generator_1.h_count[4] ),
    .A2(_1131_),
    .ZN(_1456_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3873_ (.A1(_1268_),
    .A2(_1456_),
    .ZN(_1457_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _3874_ (.A1(_1132_),
    .A2(_1249_),
    .A3(_1455_),
    .A4(_1457_),
    .ZN(_1458_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _3875_ (.A1(net18),
    .A2(_1458_),
    .Z(_1459_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3876_ (.I(_1459_),
    .Z(_1460_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3877_ (.A1(_1216_),
    .A2(_1460_),
    .ZN(_0013_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3878_ (.I(_0689_),
    .Z(_1461_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _3879_ (.A1(_1461_),
    .A2(_1268_),
    .A3(_1281_),
    .ZN(_0014_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3880_ (.I(_1460_),
    .ZN(_1462_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3881_ (.A1(\soc.video_generator_1.h_count[2] ),
    .A2(_1281_),
    .B(_1462_),
    .ZN(_1463_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3882_ (.A1(\soc.video_generator_1.h_count[2] ),
    .A2(_1281_),
    .B(_1463_),
    .ZN(_0015_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _3883_ (.A1(\soc.video_generator_1.h_count[3] ),
    .A2(\soc.video_generator_1.h_count[2] ),
    .A3(_1281_),
    .Z(_1464_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3884_ (.A1(\soc.video_generator_1.h_count[2] ),
    .A2(_1281_),
    .B(\soc.video_generator_1.h_count[3] ),
    .ZN(_1465_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _3885_ (.A1(_1460_),
    .A2(_1464_),
    .A3(_1465_),
    .ZN(_0016_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3886_ (.A1(\soc.video_generator_1.h_count[4] ),
    .A2(_1464_),
    .Z(_1466_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3887_ (.A1(\soc.video_generator_1.h_count[4] ),
    .A2(_1464_),
    .ZN(_1467_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _3888_ (.A1(_1460_),
    .A2(_1466_),
    .A3(_1467_),
    .ZN(_0017_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3889_ (.A1(_1190_),
    .A2(_1466_),
    .B(_1462_),
    .ZN(_1468_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3890_ (.A1(_1190_),
    .A2(_1466_),
    .B(_1468_),
    .ZN(_0018_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3891_ (.A1(_1190_),
    .A2(_1466_),
    .B(_1131_),
    .ZN(_1469_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _3892_ (.A1(_1190_),
    .A2(_1131_),
    .A3(_1466_),
    .Z(_1470_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _3893_ (.A1(_1460_),
    .A2(_1469_),
    .A3(_1470_),
    .ZN(_0019_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3894_ (.A1(_1132_),
    .A2(_1470_),
    .B(_1462_),
    .ZN(_1471_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3895_ (.A1(_1132_),
    .A2(_1470_),
    .B(_1471_),
    .ZN(_0020_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3896_ (.A1(_1132_),
    .A2(_1470_),
    .ZN(_1472_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3897_ (.A1(_1132_),
    .A2(\soc.video_generator_1.h_count[8] ),
    .A3(_1470_),
    .ZN(_1473_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3898_ (.A1(_1462_),
    .A2(_1473_),
    .ZN(_1474_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3899_ (.A1(_1130_),
    .A2(_1472_),
    .B(_1474_),
    .ZN(_0021_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3900_ (.A1(\soc.video_generator_1.h_count[9] ),
    .A2(_1473_),
    .Z(_1475_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3901_ (.A1(_1460_),
    .A2(_1475_),
    .ZN(_0022_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3902_ (.A1(\soc.rom_encoder_0.initializing_step[1] ),
    .A2(_1438_),
    .B(\soc.rom_encoder_0.initializing_step[2] ),
    .ZN(_1476_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _3903_ (.A1(\soc.rom_encoder_0.initializing_step[4] ),
    .A2(\soc.rom_encoder_0.initializing_step[3] ),
    .A3(_1476_),
    .ZN(_1477_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3904_ (.A1(_1407_),
    .A2(\soc.rom_encoder_0.current_state[1] ),
    .ZN(_1478_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3905_ (.A1(_1419_),
    .A2(_1478_),
    .ZN(_1479_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _3906_ (.A1(\soc.rom_encoder_0.output_buffer[16] ),
    .A2(_1440_),
    .A3(_1479_),
    .ZN(_1480_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3907_ (.I(_1418_),
    .Z(_1481_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3908_ (.A1(_1478_),
    .A2(_1434_),
    .B(_1421_),
    .ZN(_1482_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3909_ (.I(_1479_),
    .ZN(_1483_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _3910_ (.A1(\soc.rom_encoder_0.request_data_out[12] ),
    .A2(_1481_),
    .B1(_1482_),
    .B2(\soc.rom_encoder_0.output_buffer[16] ),
    .C(_1483_),
    .ZN(_1484_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _3911_ (.A1(_1410_),
    .A2(_1439_),
    .A3(_1477_),
    .B1(_1480_),
    .B2(_1484_),
    .ZN(_1485_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _3912_ (.A1(\soc.rom_encoder_0.initializing_step[4] ),
    .A2(\soc.rom_encoder_0.initializing_step[3] ),
    .A3(_1430_),
    .B(_1432_),
    .ZN(_1486_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _3913_ (.A1(_1430_),
    .A2(_1485_),
    .B1(_1486_),
    .B2(net64),
    .ZN(_1487_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3914_ (.A1(_0676_),
    .A2(_1487_),
    .ZN(_0023_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _3915_ (.I(\soc.ram_encoder_0.current_state[0] ),
    .Z(_1488_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _3916_ (.I(\soc.ram_encoder_0.current_state[2] ),
    .ZN(_1489_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _3917_ (.I(\soc.ram_encoder_0.current_state[1] ),
    .ZN(_1490_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _3918_ (.A1(_1489_),
    .A2(_1490_),
    .ZN(_1491_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3919_ (.A1(_1488_),
    .A2(_1491_),
    .ZN(_1492_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _3920_ (.I(\soc.ram_encoder_0.current_state[2] ),
    .Z(_1493_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _3921_ (.A1(\soc.ram_encoder_0.initializing_step[4] ),
    .A2(\soc.ram_encoder_0.initializing_step[3] ),
    .A3(\soc.ram_encoder_0.initializing_step[2] ),
    .A4(\soc.ram_encoder_0.initializing_step[1] ),
    .ZN(_1494_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _3922_ (.A1(_1488_),
    .A2(_1494_),
    .ZN(_1495_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _3923_ (.A1(\soc.ram_encoder_0.current_state[1] ),
    .A2(_1488_),
    .ZN(_1496_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3924_ (.I(\soc.ram_encoder_0.output_bits_left[3] ),
    .ZN(_1497_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3925_ (.A1(\soc.ram_encoder_0.output_bits_left[2] ),
    .A2(_1497_),
    .ZN(_1498_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _3926_ (.A1(\soc.ram_encoder_0.output_bits_left[4] ),
    .A2(_1498_),
    .ZN(_1499_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3927_ (.A1(\soc.ram_encoder_0.current_state[2] ),
    .A2(_1490_),
    .ZN(_1500_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3928_ (.A1(_1488_),
    .A2(_1500_),
    .ZN(_1501_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _3929_ (.I(\soc.ram_encoder_0.current_state[0] ),
    .ZN(_1502_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3930_ (.A1(\soc.ram_encoder_0.current_state[1] ),
    .A2(_1502_),
    .ZN(_1503_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3931_ (.A1(\soc.ram_encoder_0.current_state[2] ),
    .A2(_1503_),
    .ZN(_1504_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3932_ (.A1(\soc.ram_encoder_0.request_write ),
    .A2(_1501_),
    .B(_1504_),
    .ZN(_1505_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3933_ (.A1(_1499_),
    .A2(_1505_),
    .ZN(_1506_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3934_ (.A1(\soc.ram_encoder_0.toggled_sram_sck ),
    .A2(_1506_),
    .ZN(_1507_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _3935_ (.A1(_1493_),
    .A2(_1495_),
    .B(_1496_),
    .C(_1507_),
    .ZN(_1508_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _3936_ (.A1(_0674_),
    .A2(_1492_),
    .A3(_1508_),
    .ZN(_1509_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3937_ (.I(_1509_),
    .Z(_1510_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _3938_ (.A1(\soc.ram_encoder_0.output_bits_left[4] ),
    .A2(_1498_),
    .Z(_1511_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3939_ (.A1(\soc.ram_encoder_0.current_state[1] ),
    .A2(_1502_),
    .ZN(_1512_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _3940_ (.A1(_1493_),
    .A2(_1511_),
    .A3(_1512_),
    .ZN(_1513_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3941_ (.I(_1513_),
    .Z(_1514_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _3942_ (.A1(_1491_),
    .A2(_1496_),
    .ZN(_1515_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3943_ (.A1(\soc.ram_encoder_0.initializing_step[0] ),
    .A2(_1494_),
    .ZN(_1516_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3944_ (.A1(_1500_),
    .A2(_1511_),
    .ZN(_1517_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3945_ (.A1(_1504_),
    .A2(_1517_),
    .Z(_1518_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3946_ (.A1(_1515_),
    .A2(_1516_),
    .B(_1518_),
    .ZN(_1519_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3947_ (.I(_1519_),
    .Z(_1520_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3948_ (.A1(\soc.ram_encoder_0.request_address[4] ),
    .A2(_1514_),
    .B1(_1520_),
    .B2(\soc.ram_encoder_0.output_buffer[1] ),
    .ZN(_1521_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3949_ (.I(_1509_),
    .Z(_1522_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3950_ (.A1(\soc.ram_encoder_0.output_buffer[5] ),
    .A2(_1522_),
    .ZN(_1523_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3951_ (.A1(_1510_),
    .A2(_1521_),
    .B(_1523_),
    .ZN(_0024_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3952_ (.A1(\soc.ram_encoder_0.request_address[5] ),
    .A2(_1514_),
    .B1(_1520_),
    .B2(\soc.ram_encoder_0.output_buffer[2] ),
    .ZN(_1524_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3953_ (.A1(\soc.ram_encoder_0.output_buffer[6] ),
    .A2(_1522_),
    .ZN(_1525_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3954_ (.A1(_1510_),
    .A2(_1524_),
    .B(_1525_),
    .ZN(_0025_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3955_ (.A1(\soc.ram_encoder_0.request_address[6] ),
    .A2(_1514_),
    .B1(_1520_),
    .B2(\soc.ram_encoder_0.output_buffer[3] ),
    .ZN(_1526_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3956_ (.I(_1509_),
    .Z(_1527_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3957_ (.A1(\soc.ram_encoder_0.output_buffer[7] ),
    .A2(_1527_),
    .ZN(_1528_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3958_ (.A1(_1510_),
    .A2(_1526_),
    .B(_1528_),
    .ZN(_0026_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _3959_ (.A1(_1501_),
    .A2(_1511_),
    .ZN(_1529_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _3960_ (.I(_1529_),
    .Z(_1530_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3961_ (.A1(\soc.ram_encoder_0.request_address[7] ),
    .A2(_1514_),
    .Z(_1531_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _3962_ (.A1(\soc.ram_encoder_0.output_buffer[4] ),
    .A2(_1520_),
    .B1(_1530_),
    .B2(\soc.ram_encoder_0.request_data_out[0] ),
    .C(_1531_),
    .ZN(_1532_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3963_ (.A1(\soc.ram_encoder_0.output_buffer[8] ),
    .A2(_1527_),
    .ZN(_1533_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3964_ (.A1(_1510_),
    .A2(_1532_),
    .B(_1533_),
    .ZN(_0027_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3965_ (.A1(\soc.ram_encoder_0.request_address[8] ),
    .A2(_1513_),
    .Z(_1534_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _3966_ (.A1(\soc.ram_encoder_0.output_buffer[5] ),
    .A2(_1520_),
    .B1(_1530_),
    .B2(\soc.ram_encoder_0.request_data_out[1] ),
    .C(_1534_),
    .ZN(_1535_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3967_ (.A1(\soc.ram_encoder_0.output_buffer[9] ),
    .A2(_1527_),
    .ZN(_1536_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3968_ (.A1(_1510_),
    .A2(_1535_),
    .B(_1536_),
    .ZN(_0028_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3969_ (.A1(\soc.ram_encoder_0.request_address[9] ),
    .A2(_1513_),
    .Z(_1537_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _3970_ (.A1(\soc.ram_encoder_0.output_buffer[6] ),
    .A2(_1520_),
    .B1(_1530_),
    .B2(\soc.ram_encoder_0.request_data_out[2] ),
    .C(_1537_),
    .ZN(_1538_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3971_ (.A1(\soc.ram_encoder_0.output_buffer[10] ),
    .A2(_1527_),
    .ZN(_1539_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3972_ (.A1(_1510_),
    .A2(_1538_),
    .B(_1539_),
    .ZN(_0029_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3973_ (.A1(\soc.ram_encoder_0.request_address[10] ),
    .A2(_1513_),
    .Z(_1540_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _3974_ (.A1(\soc.ram_encoder_0.output_buffer[7] ),
    .A2(_1520_),
    .B1(_1530_),
    .B2(\soc.ram_encoder_0.request_data_out[3] ),
    .C(_1540_),
    .ZN(_1541_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3975_ (.A1(\soc.ram_encoder_0.output_buffer[11] ),
    .A2(_1527_),
    .ZN(_1542_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3976_ (.A1(_1510_),
    .A2(_1541_),
    .B(_1542_),
    .ZN(_0030_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3977_ (.A1(\soc.ram_encoder_0.request_address[11] ),
    .A2(_1513_),
    .Z(_1543_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _3978_ (.A1(\soc.ram_encoder_0.output_buffer[8] ),
    .A2(_1520_),
    .B1(_1530_),
    .B2(\soc.ram_encoder_0.request_data_out[4] ),
    .C(_1543_),
    .ZN(_1544_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3979_ (.A1(\soc.ram_encoder_0.output_buffer[12] ),
    .A2(_1527_),
    .ZN(_1545_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3980_ (.A1(_1510_),
    .A2(_1544_),
    .B(_1545_),
    .ZN(_0031_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3981_ (.A1(\soc.ram_encoder_0.request_address[12] ),
    .A2(_1513_),
    .Z(_1546_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _3982_ (.A1(\soc.ram_encoder_0.output_buffer[9] ),
    .A2(_1520_),
    .B1(_1530_),
    .B2(\soc.ram_encoder_0.request_data_out[5] ),
    .C(_1546_),
    .ZN(_1547_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3983_ (.A1(\soc.ram_encoder_0.output_buffer[13] ),
    .A2(_1527_),
    .ZN(_1548_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3984_ (.A1(_1510_),
    .A2(_1547_),
    .B(_1548_),
    .ZN(_0032_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3985_ (.A1(\soc.ram_encoder_0.request_address[13] ),
    .A2(_1513_),
    .Z(_1549_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _3986_ (.A1(\soc.ram_encoder_0.output_buffer[10] ),
    .A2(_1520_),
    .B1(_1530_),
    .B2(\soc.ram_encoder_0.request_data_out[6] ),
    .C(_1549_),
    .ZN(_1550_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3987_ (.A1(\soc.ram_encoder_0.output_buffer[14] ),
    .A2(_1527_),
    .ZN(_1551_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3988_ (.A1(_1510_),
    .A2(_1550_),
    .B(_1551_),
    .ZN(_0033_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3989_ (.A1(\soc.ram_encoder_0.output_buffer[11] ),
    .A2(_1519_),
    .Z(_1552_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _3990_ (.A1(\soc.ram_encoder_0.request_address[14] ),
    .A2(_1514_),
    .B1(_1530_),
    .B2(\soc.ram_encoder_0.request_data_out[7] ),
    .C(_1552_),
    .ZN(_1553_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3991_ (.A1(\soc.ram_encoder_0.output_buffer[15] ),
    .A2(_1527_),
    .ZN(_1554_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3992_ (.A1(_1522_),
    .A2(_1553_),
    .B(_1554_),
    .ZN(_0034_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3993_ (.A1(_1515_),
    .A2(_1518_),
    .ZN(_1555_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3994_ (.A1(\soc.ram_encoder_0.output_buffer[12] ),
    .A2(_1555_),
    .ZN(_1556_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _3995_ (.A1(_1493_),
    .A2(\soc.ram_encoder_0.current_state[1] ),
    .A3(_1502_),
    .ZN(_1557_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3996_ (.I(\soc.ram_encoder_0.request_write ),
    .ZN(_1558_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _3997_ (.A1(\soc.ram_encoder_0.initializing_step[0] ),
    .A2(_1494_),
    .B(_1515_),
    .ZN(_1559_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _3998_ (.A1(\soc.ram_encoder_0.request_data_out[8] ),
    .A2(_1529_),
    .B1(_1557_),
    .B2(_1558_),
    .C(_1559_),
    .ZN(_1560_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3999_ (.A1(_1556_),
    .A2(_1560_),
    .ZN(_1561_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4000_ (.I0(_1561_),
    .I1(\soc.ram_encoder_0.output_buffer[16] ),
    .S(_1509_),
    .Z(_1562_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4001_ (.I(_1562_),
    .Z(_0035_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4002_ (.A1(\soc.ram_encoder_0.request_data_out[9] ),
    .A2(_1515_),
    .A3(_1529_),
    .ZN(_1563_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4003_ (.A1(_1499_),
    .A2(_1515_),
    .ZN(_1564_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4004_ (.A1(\soc.ram_encoder_0.output_buffer[13] ),
    .A2(_1564_),
    .ZN(_1565_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4005_ (.A1(_1563_),
    .A2(_1565_),
    .ZN(_1566_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _4006_ (.A1(_1557_),
    .A2(_1559_),
    .A3(_1566_),
    .ZN(_1567_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4007_ (.A1(\soc.ram_encoder_0.output_buffer[17] ),
    .A2(_1527_),
    .ZN(_1568_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4008_ (.A1(_1522_),
    .A2(_1567_),
    .B(_1568_),
    .ZN(_0036_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _4009_ (.A1(\soc.ram_encoder_0.output_buffer[14] ),
    .A2(_1555_),
    .B1(_1530_),
    .B2(\soc.ram_encoder_0.request_data_out[10] ),
    .C(_1559_),
    .ZN(_1569_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4010_ (.A1(\soc.ram_encoder_0.output_buffer[18] ),
    .A2(_1509_),
    .ZN(_1570_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4011_ (.A1(_1522_),
    .A2(_1569_),
    .B(_1570_),
    .ZN(_0037_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _4012_ (.A1(\soc.ram_encoder_0.output_buffer[15] ),
    .A2(_1555_),
    .B1(_1530_),
    .B2(\soc.ram_encoder_0.request_data_out[11] ),
    .C(_1559_),
    .ZN(_1571_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4013_ (.A1(\soc.ram_encoder_0.output_buffer[19] ),
    .A2(_1509_),
    .ZN(_1572_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4014_ (.A1(_1522_),
    .A2(_1571_),
    .B(_1572_),
    .ZN(_0038_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4015_ (.A1(\soc.spi_video_ram_1.current_state[3] ),
    .A2(\soc.spi_video_ram_1.current_state[0] ),
    .ZN(_1573_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4016_ (.A1(\soc.spi_video_ram_1.current_state[4] ),
    .A2(_0725_),
    .B(_0685_),
    .ZN(_1574_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4017_ (.A1(\soc.spi_video_ram_1.state_sram_clk_counter[1] ),
    .A2(_0685_),
    .ZN(_1575_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _4018_ (.A1(_1573_),
    .A2(_1574_),
    .B(_1575_),
    .ZN(_1576_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4019_ (.A1(_0674_),
    .A2(_0706_),
    .ZN(_0188_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4020_ (.A1(_1576_),
    .A2(_0188_),
    .Z(_1577_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _4021_ (.I(_1577_),
    .Z(_1578_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4022_ (.I(_0002_),
    .Z(_1579_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4023_ (.I(_1579_),
    .Z(_1580_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4024_ (.I(_1580_),
    .Z(_1581_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 _4025_ (.I(_0000_),
    .Z(_1582_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _4026_ (.I(_1582_),
    .Z(_1583_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 _4027_ (.I(_1583_),
    .Z(_1584_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 _4028_ (.I(_1584_),
    .Z(_1585_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4029_ (.I(_0001_),
    .Z(_1586_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _4030_ (.I(_1586_),
    .Z(_1587_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4031_ (.I(_1587_),
    .Z(_1588_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4032_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[0][16] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[1][16] ),
    .I2(\soc.spi_video_ram_1.write_fifo.fifo_mem[2][16] ),
    .I3(\soc.spi_video_ram_1.write_fifo.fifo_mem[3][16] ),
    .S0(_1585_),
    .S1(_1588_),
    .Z(_1589_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4033_ (.I(_0001_),
    .Z(_1590_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4034_ (.I(_1590_),
    .Z(_1591_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4035_ (.I(_1591_),
    .Z(_1592_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 _4036_ (.I(_1583_),
    .Z(_1593_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 _4037_ (.I(_1593_),
    .Z(_1594_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4038_ (.I(_1594_),
    .Z(_1595_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4039_ (.I(_1584_),
    .Z(_1596_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4040_ (.I(\soc.spi_video_ram_1.write_fifo.fifo_mem[5][16] ),
    .ZN(_1597_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4041_ (.A1(_1596_),
    .A2(_1597_),
    .ZN(_1598_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4042_ (.A1(_1595_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[4][16] ),
    .B(_1598_),
    .ZN(_1599_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 _4043_ (.I(_1583_),
    .Z(_1600_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4044_ (.I(_1600_),
    .Z(_1601_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4045_ (.I(\soc.spi_video_ram_1.write_fifo.fifo_mem[7][16] ),
    .ZN(_1602_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4046_ (.A1(_1594_),
    .A2(_1602_),
    .ZN(_1603_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4047_ (.A1(_1601_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[6][16] ),
    .B(_1603_),
    .C(_1588_),
    .ZN(_1604_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4048_ (.I(_1579_),
    .Z(_1605_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4049_ (.A1(_1592_),
    .A2(_1599_),
    .B(_1604_),
    .C(_1605_),
    .ZN(_1606_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _4050_ (.A1(\soc.spi_video_ram_1.state_sram_clk_counter[8] ),
    .A2(\soc.spi_video_ram_1.state_sram_clk_counter[0] ),
    .A3(_0684_),
    .ZN(_1607_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4051_ (.A1(\soc.spi_video_ram_1.state_sram_clk_counter[1] ),
    .A2(_1607_),
    .ZN(_1608_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _4052_ (.A1(_0710_),
    .A2(_1608_),
    .ZN(_1609_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4053_ (.A1(_1581_),
    .A2(_1589_),
    .B(_1606_),
    .C(_1609_),
    .ZN(_1610_));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _4054_ (.A1(_0689_),
    .A2(_0705_),
    .A3(_1576_),
    .Z(_1611_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4055_ (.I(_1611_),
    .Z(_1612_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4056_ (.A1(\soc.spi_video_ram_1.output_buffer[1] ),
    .A2(_1612_),
    .ZN(_1613_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4057_ (.A1(_1578_),
    .A2(_1610_),
    .B(_1613_),
    .ZN(_0039_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4058_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[0][18] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[1][18] ),
    .I2(\soc.spi_video_ram_1.write_fifo.fifo_mem[2][18] ),
    .I3(\soc.spi_video_ram_1.write_fifo.fifo_mem[3][18] ),
    .S0(_1585_),
    .S1(_1588_),
    .Z(_1614_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4059_ (.I(\soc.spi_video_ram_1.write_fifo.fifo_mem[5][18] ),
    .ZN(_1615_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4060_ (.A1(_1596_),
    .A2(_1615_),
    .ZN(_1616_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4061_ (.A1(_1595_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[4][18] ),
    .B(_1616_),
    .ZN(_1617_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4062_ (.I(\soc.spi_video_ram_1.write_fifo.fifo_mem[7][18] ),
    .ZN(_1618_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4063_ (.A1(_1594_),
    .A2(_1618_),
    .ZN(_1619_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4064_ (.A1(_1601_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[6][18] ),
    .B(_1619_),
    .C(_1588_),
    .ZN(_1620_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4065_ (.A1(_1592_),
    .A2(_1617_),
    .B(_1620_),
    .C(_1605_),
    .ZN(_1621_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4066_ (.A1(_1581_),
    .A2(_1614_),
    .B(_1621_),
    .C(_1609_),
    .ZN(_1622_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4067_ (.A1(\soc.spi_video_ram_1.output_buffer[3] ),
    .A2(_1612_),
    .ZN(_1623_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4068_ (.A1(_1578_),
    .A2(_1622_),
    .B(_1623_),
    .ZN(_0040_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4069_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[0][17] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[1][17] ),
    .I2(\soc.spi_video_ram_1.write_fifo.fifo_mem[2][17] ),
    .I3(\soc.spi_video_ram_1.write_fifo.fifo_mem[3][17] ),
    .S0(_1585_),
    .S1(_1588_),
    .Z(_1624_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4070_ (.I(\soc.spi_video_ram_1.write_fifo.fifo_mem[5][17] ),
    .ZN(_1625_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4071_ (.A1(_1596_),
    .A2(_1625_),
    .ZN(_1626_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4072_ (.A1(_1601_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[4][17] ),
    .B(_1626_),
    .ZN(_1627_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4073_ (.I(\soc.spi_video_ram_1.write_fifo.fifo_mem[7][17] ),
    .ZN(_1628_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4074_ (.A1(_1594_),
    .A2(_1628_),
    .ZN(_1629_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4075_ (.A1(_1601_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[6][17] ),
    .B(_1629_),
    .C(_1591_),
    .ZN(_1630_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4076_ (.A1(_1592_),
    .A2(_1627_),
    .B(_1630_),
    .C(_1605_),
    .ZN(_1631_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4077_ (.A1(_1581_),
    .A2(_1624_),
    .B(_1631_),
    .C(_1609_),
    .ZN(_1632_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4078_ (.A1(\soc.spi_video_ram_1.output_buffer[2] ),
    .A2(_1612_),
    .ZN(_1633_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4079_ (.A1(_1578_),
    .A2(_1632_),
    .B(_1633_),
    .ZN(_0041_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _4080_ (.A1(_0674_),
    .A2(\soc.ram_encoder_0.toggled_sram_sck ),
    .A3(_1506_),
    .A4(_1515_),
    .ZN(_1634_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4081_ (.I(_1634_),
    .ZN(_1635_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4082_ (.A1(_1497_),
    .A2(\soc.ram_encoder_0.output_bits_left[4] ),
    .ZN(_1636_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4083_ (.A1(_1493_),
    .A2(_1490_),
    .B(_1504_),
    .ZN(_1637_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4084_ (.A1(\soc.ram_encoder_0.output_bits_left[2] ),
    .A2(_1636_),
    .B(_1637_),
    .ZN(_1638_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4085_ (.A1(_1497_),
    .A2(_1635_),
    .B(\soc.ram_encoder_0.output_bits_left[4] ),
    .ZN(_1639_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4086_ (.A1(_1635_),
    .A2(_1638_),
    .B(_1639_),
    .ZN(_0042_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4087_ (.A1(\soc.ram_encoder_0.output_bits_left[2] ),
    .A2(\soc.ram_encoder_0.output_bits_left[3] ),
    .Z(_1640_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4088_ (.A1(_1637_),
    .A2(_1640_),
    .ZN(_1641_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _4089_ (.A1(_1514_),
    .A2(_1634_),
    .A3(_1641_),
    .ZN(_1642_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4090_ (.A1(_1497_),
    .A2(_1634_),
    .B(_1642_),
    .ZN(_0043_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _4091_ (.A1(\soc.ram_encoder_0.output_bits_left[2] ),
    .A2(_1557_),
    .A3(_1634_),
    .Z(_1643_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4092_ (.A1(\soc.ram_encoder_0.output_bits_left[2] ),
    .A2(_1634_),
    .ZN(_1644_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4093_ (.A1(_1643_),
    .A2(_1644_),
    .ZN(_0044_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _4094_ (.A1(_0674_),
    .A2(_1427_),
    .A3(_1424_),
    .ZN(_1645_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4095_ (.I(_1645_),
    .ZN(_1646_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4096_ (.A1(_1415_),
    .A2(_1646_),
    .ZN(_1647_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4097_ (.A1(_1478_),
    .A2(_1421_),
    .ZN(_1648_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _4098_ (.A1(\soc.rom_encoder_0.output_bits_left[2] ),
    .A2(_1414_),
    .A3(\soc.rom_encoder_0.output_bits_left[3] ),
    .B(_1648_),
    .ZN(_1649_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4099_ (.A1(_1414_),
    .A2(_1647_),
    .B1(_1649_),
    .B2(_1646_),
    .ZN(_0045_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _4100_ (.A1(_1406_),
    .A2(_1478_),
    .A3(_1417_),
    .ZN(_1650_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4101_ (.I(_1650_),
    .ZN(_1651_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4102_ (.I(\soc.rom_encoder_0.output_bits_left[2] ),
    .ZN(_1652_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4103_ (.A1(_1652_),
    .A2(\soc.rom_encoder_0.output_bits_left[3] ),
    .ZN(_1653_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4104_ (.A1(_1433_),
    .A2(_1653_),
    .ZN(_1654_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _4105_ (.A1(_1646_),
    .A2(_1648_),
    .A3(_1651_),
    .A4(_1654_),
    .Z(_1655_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4106_ (.A1(_1415_),
    .A2(_1645_),
    .B(_1655_),
    .ZN(_0046_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4107_ (.A1(_1408_),
    .A2(_1435_),
    .ZN(_1656_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4108_ (.A1(_1652_),
    .A2(_1656_),
    .B(_1645_),
    .ZN(_1657_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4109_ (.A1(_1652_),
    .A2(_1645_),
    .B(_1657_),
    .ZN(_0047_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4110_ (.I(\soc.cpu.AReg.data[15] ),
    .ZN(_1658_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4111_ (.A1(_1111_),
    .A2(_1114_),
    .ZN(_1659_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4112_ (.A1(_0954_),
    .A2(_1659_),
    .ZN(_1660_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4113_ (.A1(_1120_),
    .A2(_1660_),
    .Z(_1661_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4114_ (.A1(_0907_),
    .A2(\soc.cpu.AReg.data[15] ),
    .B1(_1012_),
    .B2(\soc.ram_data_out[15] ),
    .ZN(_1662_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4115_ (.A1(_1011_),
    .A2(_1662_),
    .ZN(_1663_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4116_ (.A1(_0926_),
    .A2(_1663_),
    .ZN(_1664_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4117_ (.A1(_0904_),
    .A2(\soc.cpu.ALU.x[15] ),
    .ZN(_1665_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4118_ (.A1(_0923_),
    .A2(_1665_),
    .ZN(_1666_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4119_ (.A1(_0954_),
    .A2(_1664_),
    .B(_1666_),
    .ZN(_1667_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4120_ (.A1(_1664_),
    .A2(_1666_),
    .B(_1667_),
    .ZN(_1668_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _4121_ (.A1(_0990_),
    .A2(_1661_),
    .A3(_1668_),
    .Z(_1669_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _4122_ (.A1(_1658_),
    .A2(_0881_),
    .B1(_1669_),
    .B2(_0848_),
    .ZN(_0048_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _4123_ (.A1(_0674_),
    .A2(_1410_),
    .A3(_1431_),
    .ZN(_1670_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4124_ (.I(_1670_),
    .Z(_1671_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4125_ (.A1(_1651_),
    .A2(_1670_),
    .ZN(_1672_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4126_ (.A1(\soc.rom_encoder_0.output_buffer[4] ),
    .A2(_1671_),
    .B1(_1672_),
    .B2(\soc.rom_encoder_0.request_address[3] ),
    .ZN(_1673_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4127_ (.I(_1673_),
    .ZN(_0049_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4128_ (.A1(\soc.rom_encoder_0.output_buffer[3] ),
    .A2(_1671_),
    .B1(_1672_),
    .B2(\soc.rom_encoder_0.request_address[2] ),
    .ZN(_1674_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4129_ (.I(_1674_),
    .ZN(_0050_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4130_ (.A1(\soc.rom_encoder_0.output_buffer[2] ),
    .A2(_1671_),
    .B1(_1672_),
    .B2(\soc.rom_encoder_0.request_address[1] ),
    .ZN(_1675_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4131_ (.I(_1675_),
    .ZN(_0051_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4132_ (.A1(\soc.rom_encoder_0.output_buffer[1] ),
    .A2(_1671_),
    .B1(_1672_),
    .B2(\soc.rom_encoder_0.request_address[0] ),
    .ZN(_1676_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4133_ (.I(_1676_),
    .ZN(_0052_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4134_ (.A1(\soc.ram_encoder_0.request_address[3] ),
    .A2(_1514_),
    .ZN(_1677_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4135_ (.A1(\soc.ram_encoder_0.output_buffer[4] ),
    .A2(_1509_),
    .ZN(_1678_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4136_ (.A1(_1522_),
    .A2(_1677_),
    .B(_1678_),
    .ZN(_0053_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4137_ (.A1(\soc.ram_encoder_0.request_address[2] ),
    .A2(_1514_),
    .ZN(_1679_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4138_ (.A1(\soc.ram_encoder_0.output_buffer[3] ),
    .A2(_1509_),
    .ZN(_1680_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4139_ (.A1(_1522_),
    .A2(_1679_),
    .B(_1680_),
    .ZN(_0054_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4140_ (.A1(\soc.ram_encoder_0.request_address[1] ),
    .A2(_1514_),
    .ZN(_1681_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4141_ (.A1(\soc.ram_encoder_0.output_buffer[2] ),
    .A2(_1509_),
    .ZN(_1682_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4142_ (.A1(_1522_),
    .A2(_1681_),
    .B(_1682_),
    .ZN(_0055_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4143_ (.A1(\soc.ram_encoder_0.request_address[0] ),
    .A2(_1514_),
    .ZN(_1683_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4144_ (.A1(\soc.ram_encoder_0.output_buffer[1] ),
    .A2(_1509_),
    .ZN(_1684_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4145_ (.A1(_1522_),
    .A2(_1683_),
    .B(_1684_),
    .ZN(_0056_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4146_ (.I(\soc.spi_video_ram_1.output_buffer[23] ),
    .ZN(_1685_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4147_ (.I(_1611_),
    .Z(_1686_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4148_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[0][0] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[1][0] ),
    .I2(\soc.spi_video_ram_1.write_fifo.fifo_mem[2][0] ),
    .I3(\soc.spi_video_ram_1.write_fifo.fifo_mem[3][0] ),
    .S0(_1594_),
    .S1(_1588_),
    .Z(_1687_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4149_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[4][0] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[5][0] ),
    .I2(\soc.spi_video_ram_1.write_fifo.fifo_mem[6][0] ),
    .I3(\soc.spi_video_ram_1.write_fifo.fifo_mem[7][0] ),
    .S0(_1593_),
    .S1(_1587_),
    .Z(_1688_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4150_ (.I(_1688_),
    .ZN(_1689_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4151_ (.A1(_1605_),
    .A2(_1689_),
    .ZN(_1690_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4152_ (.A1(_1581_),
    .A2(_1687_),
    .B(_1690_),
    .C(_0685_),
    .ZN(_1691_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4153_ (.A1(_0720_),
    .A2(_0704_),
    .ZN(_1692_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _4154_ (.A1(_1352_),
    .A2(_1353_),
    .A3(_1354_),
    .ZN(_1693_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4155_ (.A1(_0681_),
    .A2(_1607_),
    .ZN(_1694_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4156_ (.A1(\soc.spi_video_ram_1.current_state[4] ),
    .A2(_1694_),
    .ZN(_1695_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4157_ (.A1(_1693_),
    .A2(_1695_),
    .ZN(_1696_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _4158_ (.A1(_1692_),
    .A2(_1578_),
    .A3(_1696_),
    .ZN(_1697_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4159_ (.A1(_1685_),
    .A2(_1686_),
    .B1(_1691_),
    .B2(_1697_),
    .ZN(_0057_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4160_ (.I(\soc.spi_video_ram_1.write_fifo.fifo_mem[1][1] ),
    .ZN(_1698_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4161_ (.A1(_1601_),
    .A2(_1698_),
    .B(_1591_),
    .ZN(_1699_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4162_ (.A1(_1595_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[0][1] ),
    .B(_1699_),
    .ZN(_1700_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4163_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[2][1] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[3][1] ),
    .S(_1600_),
    .Z(_1701_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4164_ (.I(_1579_),
    .Z(_1702_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4165_ (.A1(_1592_),
    .A2(_1701_),
    .B(_1702_),
    .ZN(_1703_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4166_ (.A1(_1700_),
    .A2(_1703_),
    .ZN(_1704_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4167_ (.I(\soc.spi_video_ram_1.write_fifo.fifo_mem[5][1] ),
    .ZN(_1705_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4168_ (.A1(_1596_),
    .A2(_1705_),
    .ZN(_1706_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4169_ (.A1(_1595_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[4][1] ),
    .B(_1706_),
    .ZN(_1707_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4170_ (.I(\soc.spi_video_ram_1.write_fifo.fifo_mem[7][1] ),
    .ZN(_1708_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4171_ (.A1(_1585_),
    .A2(_1708_),
    .ZN(_1709_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4172_ (.I(_1586_),
    .Z(_1710_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4173_ (.I(_1710_),
    .Z(_1711_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4174_ (.A1(_1595_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[6][1] ),
    .B(_1709_),
    .C(_1711_),
    .ZN(_1712_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4175_ (.A1(_1592_),
    .A2(_1707_),
    .B(_1712_),
    .C(_1605_),
    .ZN(_1713_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4176_ (.A1(_0685_),
    .A2(_1704_),
    .A3(_1713_),
    .ZN(_1714_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4177_ (.A1(_0820_),
    .A2(_1686_),
    .B1(_1697_),
    .B2(_1714_),
    .ZN(_0058_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4178_ (.I(\soc.spi_video_ram_1.output_buffer[21] ),
    .ZN(_1715_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4179_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[0][2] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[1][2] ),
    .I2(\soc.spi_video_ram_1.write_fifo.fifo_mem[2][2] ),
    .I3(\soc.spi_video_ram_1.write_fifo.fifo_mem[3][2] ),
    .S0(_1594_),
    .S1(_1588_),
    .Z(_1716_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4180_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[4][2] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[5][2] ),
    .I2(\soc.spi_video_ram_1.write_fifo.fifo_mem[6][2] ),
    .I3(\soc.spi_video_ram_1.write_fifo.fifo_mem[7][2] ),
    .S0(_1593_),
    .S1(_1587_),
    .Z(_1717_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4181_ (.I(_1717_),
    .ZN(_1718_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4182_ (.A1(_1605_),
    .A2(_1718_),
    .ZN(_1719_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4183_ (.A1(_0710_),
    .A2(_1607_),
    .ZN(_1720_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4184_ (.A1(_1581_),
    .A2(_1716_),
    .B(_1719_),
    .C(_1720_),
    .ZN(_1721_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _4185_ (.A1(_0720_),
    .A2(_1692_),
    .A3(_1578_),
    .A4(_1696_),
    .ZN(_1722_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4186_ (.A1(_1715_),
    .A2(_1686_),
    .B1(_1721_),
    .B2(_1722_),
    .ZN(_0059_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4187_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[0][3] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[1][3] ),
    .I2(\soc.spi_video_ram_1.write_fifo.fifo_mem[2][3] ),
    .I3(\soc.spi_video_ram_1.write_fifo.fifo_mem[3][3] ),
    .S0(_1585_),
    .S1(_1711_),
    .Z(_1723_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _4188_ (.I(_1583_),
    .Z(_1724_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4189_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[4][3] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[5][3] ),
    .I2(\soc.spi_video_ram_1.write_fifo.fifo_mem[6][3] ),
    .I3(\soc.spi_video_ram_1.write_fifo.fifo_mem[7][3] ),
    .S0(_1724_),
    .S1(_1587_),
    .Z(_1725_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4190_ (.I(_1725_),
    .ZN(_1726_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4191_ (.A1(_1581_),
    .A2(_1726_),
    .ZN(_1727_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4192_ (.A1(_1581_),
    .A2(_1723_),
    .B(_1727_),
    .C(_1720_),
    .ZN(_1728_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4193_ (.A1(_0828_),
    .A2(_1686_),
    .B1(_1722_),
    .B2(_1728_),
    .ZN(_0060_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4194_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[0][4] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[1][4] ),
    .I2(\soc.spi_video_ram_1.write_fifo.fifo_mem[2][4] ),
    .I3(\soc.spi_video_ram_1.write_fifo.fifo_mem[3][4] ),
    .S0(_1585_),
    .S1(_1711_),
    .Z(_1729_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4195_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[4][4] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[5][4] ),
    .I2(\soc.spi_video_ram_1.write_fifo.fifo_mem[6][4] ),
    .I3(\soc.spi_video_ram_1.write_fifo.fifo_mem[7][4] ),
    .S0(_1593_),
    .S1(_1587_),
    .Z(_1730_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4196_ (.I(_1730_),
    .ZN(_1731_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4197_ (.A1(_1605_),
    .A2(_1731_),
    .ZN(_1732_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4198_ (.A1(_1581_),
    .A2(_1729_),
    .B(_1732_),
    .C(_1720_),
    .ZN(_1733_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4199_ (.A1(_0800_),
    .A2(_1686_),
    .B1(_1722_),
    .B2(_1733_),
    .ZN(_0061_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4200_ (.I(\soc.spi_video_ram_1.write_fifo.fifo_mem[1][5] ),
    .ZN(_1734_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4201_ (.A1(_1601_),
    .A2(_1734_),
    .B(_1591_),
    .ZN(_1735_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4202_ (.A1(_1595_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[0][5] ),
    .B(_1735_),
    .ZN(_1736_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4203_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[2][5] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[3][5] ),
    .S(_1600_),
    .Z(_1737_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4204_ (.A1(_1711_),
    .A2(_1737_),
    .B(_1702_),
    .ZN(_1738_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4205_ (.A1(_1736_),
    .A2(_1738_),
    .ZN(_1739_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4206_ (.I(\soc.spi_video_ram_1.write_fifo.fifo_mem[5][5] ),
    .ZN(_1740_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4207_ (.A1(_1596_),
    .A2(_1740_),
    .ZN(_1741_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4208_ (.A1(_1595_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[4][5] ),
    .B(_1741_),
    .ZN(_1742_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4209_ (.I(\soc.spi_video_ram_1.write_fifo.fifo_mem[7][5] ),
    .ZN(_1743_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4210_ (.A1(_1585_),
    .A2(_1743_),
    .ZN(_1744_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4211_ (.A1(_1595_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[6][5] ),
    .B(_1744_),
    .C(_1711_),
    .ZN(_1745_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4212_ (.A1(_1592_),
    .A2(_1742_),
    .B(_1745_),
    .C(_1605_),
    .ZN(_1746_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4213_ (.A1(_0685_),
    .A2(_1739_),
    .A3(_1746_),
    .ZN(_1747_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4214_ (.A1(_0801_),
    .A2(_1686_),
    .B1(_1697_),
    .B2(_1747_),
    .ZN(_0062_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4215_ (.I(\soc.spi_video_ram_1.write_fifo.fifo_mem[3][6] ),
    .ZN(_1748_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4216_ (.A1(_1594_),
    .A2(_1748_),
    .ZN(_1749_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4217_ (.A1(_1601_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[2][6] ),
    .B(_1749_),
    .ZN(_1750_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4218_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[0][6] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[1][6] ),
    .S(_1724_),
    .Z(_1751_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4219_ (.A1(_1588_),
    .A2(_1751_),
    .ZN(_1752_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _4220_ (.A1(_1592_),
    .A2(_1750_),
    .B(_1752_),
    .C(_1605_),
    .ZN(_1753_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4221_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[4][6] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[5][6] ),
    .S(_1600_),
    .Z(_1754_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _4222_ (.I(_1582_),
    .Z(_1755_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4223_ (.I(_1755_),
    .Z(_1756_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4224_ (.I(\soc.spi_video_ram_1.write_fifo.fifo_mem[7][6] ),
    .ZN(_1757_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4225_ (.A1(_1724_),
    .A2(_1757_),
    .ZN(_1758_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4226_ (.A1(_1756_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[6][6] ),
    .B(_1758_),
    .ZN(_1759_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4227_ (.A1(_1591_),
    .A2(_1759_),
    .ZN(_1760_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4228_ (.I(_1579_),
    .Z(_1761_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4229_ (.A1(_1711_),
    .A2(_1754_),
    .B(_1760_),
    .C(_1761_),
    .ZN(_1762_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4230_ (.A1(_0685_),
    .A2(_1762_),
    .ZN(_1763_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4231_ (.A1(_1753_),
    .A2(_1763_),
    .B(_0703_),
    .C(_1608_),
    .ZN(_1764_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4232_ (.A1(_1693_),
    .A2(_1694_),
    .ZN(_1765_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _4233_ (.A1(_0729_),
    .A2(_1765_),
    .B(_1578_),
    .C(_1692_),
    .ZN(_1766_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4234_ (.A1(_0799_),
    .A2(_1686_),
    .B1(_1764_),
    .B2(_1766_),
    .ZN(_0063_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4235_ (.I(\soc.spi_video_ram_1.write_fifo.fifo_mem[5][7] ),
    .ZN(_1767_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4236_ (.A1(_1601_),
    .A2(_1767_),
    .ZN(_1768_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4237_ (.A1(_1595_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[4][7] ),
    .B(_1768_),
    .ZN(_1769_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4238_ (.I(\soc.spi_video_ram_1.write_fifo.fifo_mem[7][7] ),
    .ZN(_1770_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4239_ (.A1(_1596_),
    .A2(_1770_),
    .ZN(_1771_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4240_ (.A1(_1595_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[6][7] ),
    .B(_1771_),
    .C(_1711_),
    .ZN(_1772_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4241_ (.A1(_1592_),
    .A2(_1769_),
    .B(_1772_),
    .C(_1605_),
    .ZN(_1773_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4242_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[2][7] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[3][7] ),
    .S(_1600_),
    .Z(_1774_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4243_ (.I(\soc.spi_video_ram_1.write_fifo.fifo_mem[1][7] ),
    .ZN(_1775_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4244_ (.A1(_1756_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[0][7] ),
    .ZN(_1776_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _4245_ (.A1(_1596_),
    .A2(_1775_),
    .B(_1776_),
    .C(_1591_),
    .ZN(_1777_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _4246_ (.A1(_1711_),
    .A2(_1774_),
    .B(_1777_),
    .C(_1702_),
    .ZN(_1778_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4247_ (.A1(_1607_),
    .A2(_1778_),
    .ZN(_1779_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4248_ (.A1(_1773_),
    .A2(_1779_),
    .ZN(_1780_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4249_ (.A1(_0802_),
    .A2(_1686_),
    .B1(_1766_),
    .B2(_1780_),
    .ZN(_0064_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4250_ (.I(\soc.spi_video_ram_1.write_fifo.fifo_mem[1][8] ),
    .ZN(_1781_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4251_ (.A1(_1600_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[0][8] ),
    .ZN(_1782_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _4252_ (.A1(_1594_),
    .A2(_1781_),
    .B(_1782_),
    .C(_1710_),
    .ZN(_1783_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4253_ (.I(\soc.spi_video_ram_1.write_fifo.fifo_mem[3][8] ),
    .ZN(_1784_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4254_ (.A1(_1600_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[2][8] ),
    .B(_1587_),
    .ZN(_1785_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4255_ (.A1(_1596_),
    .A2(_1784_),
    .B(_1785_),
    .ZN(_1786_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4256_ (.I(\soc.spi_video_ram_1.write_fifo.fifo_mem[5][8] ),
    .ZN(_1787_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4257_ (.A1(_1600_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[4][8] ),
    .ZN(_1788_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _4258_ (.A1(_1585_),
    .A2(_1787_),
    .B(_1788_),
    .C(_1710_),
    .ZN(_1789_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4259_ (.I(\soc.spi_video_ram_1.write_fifo.fifo_mem[7][8] ),
    .ZN(_1790_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4260_ (.A1(_1584_),
    .A2(_1790_),
    .ZN(_1791_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4261_ (.A1(_1756_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[6][8] ),
    .B(_1791_),
    .C(_1710_),
    .ZN(_1792_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4262_ (.A1(_1580_),
    .A2(_1792_),
    .ZN(_1793_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _4263_ (.A1(_1761_),
    .A2(_1783_),
    .A3(_1786_),
    .B1(_1789_),
    .B2(_1793_),
    .ZN(_1794_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _4264_ (.A1(_1693_),
    .A2(_1695_),
    .B1(_1794_),
    .B2(_1607_),
    .ZN(_1795_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _4265_ (.A1(_0689_),
    .A2(_0705_),
    .A3(_1576_),
    .ZN(_1796_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4266_ (.I0(\soc.spi_video_ram_1.output_buffer[15] ),
    .I1(_1795_),
    .S(_1796_),
    .Z(_1797_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4267_ (.I(_1797_),
    .Z(_0065_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4268_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[2][9] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[3][9] ),
    .S(_1593_),
    .Z(_1798_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4269_ (.I(\soc.spi_video_ram_1.write_fifo.fifo_mem[1][9] ),
    .ZN(_1799_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4270_ (.A1(_1724_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[0][9] ),
    .ZN(_1800_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _4271_ (.A1(_1756_),
    .A2(_1799_),
    .B(_1800_),
    .C(_1710_),
    .ZN(_1801_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _4272_ (.A1(_1711_),
    .A2(_1798_),
    .B(_1801_),
    .C(_1761_),
    .ZN(_1802_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4273_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[6][9] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[7][9] ),
    .S(_1584_),
    .Z(_1803_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4274_ (.I(\soc.spi_video_ram_1.write_fifo.fifo_mem[5][9] ),
    .ZN(_1804_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4275_ (.A1(_1593_),
    .A2(_1804_),
    .B(_1586_),
    .ZN(_1805_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4276_ (.A1(_1756_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[4][9] ),
    .B(_1805_),
    .ZN(_1806_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4277_ (.A1(_1580_),
    .A2(_1806_),
    .ZN(_1807_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4278_ (.A1(_1711_),
    .A2(_1803_),
    .B(_1807_),
    .ZN(_1808_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4279_ (.A1(_1802_),
    .A2(_1808_),
    .ZN(_1809_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4280_ (.A1(_0729_),
    .A2(_1356_),
    .B1(_1809_),
    .B2(_1608_),
    .ZN(_1810_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4281_ (.A1(_1575_),
    .A2(_1578_),
    .Z(_1811_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4282_ (.A1(\soc.spi_video_ram_1.output_buffer[14] ),
    .A2(_1612_),
    .ZN(_1812_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4283_ (.A1(_1810_),
    .A2(_1811_),
    .B(_1812_),
    .ZN(_0066_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4284_ (.A1(_1353_),
    .A2(_1354_),
    .ZN(_1813_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4285_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[0][28] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[1][28] ),
    .I2(\soc.spi_video_ram_1.write_fifo.fifo_mem[2][28] ),
    .I3(\soc.spi_video_ram_1.write_fifo.fifo_mem[3][28] ),
    .S0(_1755_),
    .S1(_1590_),
    .Z(_1814_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4286_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[4][28] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[5][28] ),
    .I2(\soc.spi_video_ram_1.write_fifo.fifo_mem[6][28] ),
    .I3(\soc.spi_video_ram_1.write_fifo.fifo_mem[7][28] ),
    .S0(_1755_),
    .S1(_1590_),
    .Z(_1815_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4287_ (.I0(_1814_),
    .I1(_1815_),
    .S(_1580_),
    .Z(_1816_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4288_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[4][10] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[5][10] ),
    .I2(\soc.spi_video_ram_1.write_fifo.fifo_mem[6][10] ),
    .I3(\soc.spi_video_ram_1.write_fifo.fifo_mem[7][10] ),
    .S0(_1755_),
    .S1(_1590_),
    .Z(_1817_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4289_ (.I(_1817_),
    .ZN(_1818_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4290_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[0][10] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[1][10] ),
    .I2(\soc.spi_video_ram_1.write_fifo.fifo_mem[2][10] ),
    .I3(\soc.spi_video_ram_1.write_fifo.fifo_mem[3][10] ),
    .S0(_1583_),
    .S1(_1586_),
    .Z(_1819_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4291_ (.A1(_1580_),
    .A2(_1819_),
    .ZN(_1820_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4292_ (.A1(_0703_),
    .A2(_1608_),
    .ZN(_1821_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _4293_ (.A1(_1702_),
    .A2(_1818_),
    .B(_1820_),
    .C(_1821_),
    .ZN(_1822_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _4294_ (.A1(_0729_),
    .A2(_1813_),
    .B1(_1816_),
    .B2(_1609_),
    .C(_1822_),
    .ZN(_1823_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4295_ (.A1(\soc.spi_video_ram_1.output_buffer[13] ),
    .A2(_1612_),
    .ZN(_1824_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4296_ (.A1(_1811_),
    .A2(_1823_),
    .B(_1824_),
    .ZN(_0067_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4297_ (.A1(_1575_),
    .A2(_1611_),
    .ZN(_1825_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4298_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[0][11] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[1][11] ),
    .I2(\soc.spi_video_ram_1.write_fifo.fifo_mem[2][11] ),
    .I3(\soc.spi_video_ram_1.write_fifo.fifo_mem[3][11] ),
    .S0(_1584_),
    .S1(_1710_),
    .Z(_1826_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4299_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[4][11] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[5][11] ),
    .I2(\soc.spi_video_ram_1.write_fifo.fifo_mem[6][11] ),
    .I3(\soc.spi_video_ram_1.write_fifo.fifo_mem[7][11] ),
    .S0(_1583_),
    .S1(_1586_),
    .Z(_1827_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4300_ (.I(_1827_),
    .ZN(_1828_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4301_ (.A1(_1761_),
    .A2(_1828_),
    .ZN(_1829_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4302_ (.A1(_1702_),
    .A2(_1826_),
    .B(_1829_),
    .ZN(_1830_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4303_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[0][27] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[1][27] ),
    .I2(\soc.spi_video_ram_1.write_fifo.fifo_mem[2][27] ),
    .I3(\soc.spi_video_ram_1.write_fifo.fifo_mem[3][27] ),
    .S0(_1583_),
    .S1(_1586_),
    .Z(_1831_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4304_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[4][27] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[5][27] ),
    .I2(\soc.spi_video_ram_1.write_fifo.fifo_mem[6][27] ),
    .I3(\soc.spi_video_ram_1.write_fifo.fifo_mem[7][27] ),
    .S0(_1583_),
    .S1(_1586_),
    .Z(_1832_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4305_ (.I0(_1831_),
    .I1(_1832_),
    .S(_1579_),
    .Z(_1833_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4306_ (.A1(_1609_),
    .A2(_1833_),
    .ZN(_1834_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4307_ (.A1(_1127_),
    .A2(_1167_),
    .ZN(_1835_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4308_ (.A1(_1257_),
    .A2(_1835_),
    .ZN(_1836_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4309_ (.A1(_0729_),
    .A2(_1354_),
    .A3(_1836_),
    .ZN(_1837_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4310_ (.A1(_1821_),
    .A2(_1830_),
    .B(_1834_),
    .C(_1837_),
    .ZN(_1838_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4311_ (.A1(\soc.spi_video_ram_1.output_buffer[12] ),
    .A2(_1612_),
    .B1(_1825_),
    .B2(_1838_),
    .ZN(_1839_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4312_ (.I(_1839_),
    .ZN(_0068_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4313_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[0][12] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[1][12] ),
    .I2(\soc.spi_video_ram_1.write_fifo.fifo_mem[2][12] ),
    .I3(\soc.spi_video_ram_1.write_fifo.fifo_mem[3][12] ),
    .S0(_1724_),
    .S1(_1587_),
    .Z(_1840_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4314_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[4][12] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[5][12] ),
    .I2(\soc.spi_video_ram_1.write_fifo.fifo_mem[6][12] ),
    .I3(\soc.spi_video_ram_1.write_fifo.fifo_mem[7][12] ),
    .S0(_1583_),
    .S1(_1586_),
    .Z(_1841_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4315_ (.I(_1841_),
    .ZN(_1842_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4316_ (.A1(_1761_),
    .A2(_1842_),
    .ZN(_1843_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4317_ (.A1(_1702_),
    .A2(_1840_),
    .B(_1843_),
    .ZN(_1844_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4318_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[0][26] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[1][26] ),
    .I2(\soc.spi_video_ram_1.write_fifo.fifo_mem[2][26] ),
    .I3(\soc.spi_video_ram_1.write_fifo.fifo_mem[3][26] ),
    .S0(_1755_),
    .S1(_1587_),
    .Z(_1845_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4319_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[4][26] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[5][26] ),
    .I2(\soc.spi_video_ram_1.write_fifo.fifo_mem[6][26] ),
    .I3(\soc.spi_video_ram_1.write_fifo.fifo_mem[7][26] ),
    .S0(_1582_),
    .S1(_1586_),
    .Z(_1846_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4320_ (.I(_1846_),
    .ZN(_1847_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4321_ (.A1(_1580_),
    .A2(_1847_),
    .ZN(_1848_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4322_ (.A1(_1702_),
    .A2(_1845_),
    .B(_1848_),
    .ZN(_1849_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4323_ (.A1(_0703_),
    .A2(_0686_),
    .ZN(_1850_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4324_ (.A1(_1127_),
    .A2(_1167_),
    .Z(_1851_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4325_ (.A1(_1129_),
    .A2(_1851_),
    .B(_0729_),
    .ZN(_1852_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _4326_ (.A1(_1821_),
    .A2(_1844_),
    .B1(_1849_),
    .B2(_1850_),
    .C(_1852_),
    .ZN(_1853_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4327_ (.A1(\soc.spi_video_ram_1.output_buffer[11] ),
    .A2(_1612_),
    .B1(_1825_),
    .B2(_1853_),
    .ZN(_1854_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4328_ (.I(_1854_),
    .ZN(_0069_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4329_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[0][25] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[1][25] ),
    .I2(\soc.spi_video_ram_1.write_fifo.fifo_mem[2][25] ),
    .I3(\soc.spi_video_ram_1.write_fifo.fifo_mem[3][25] ),
    .S0(_1755_),
    .S1(_1590_),
    .Z(_1855_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4330_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[4][25] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[5][25] ),
    .I2(\soc.spi_video_ram_1.write_fifo.fifo_mem[6][25] ),
    .I3(\soc.spi_video_ram_1.write_fifo.fifo_mem[7][25] ),
    .S0(_1582_),
    .S1(_0001_),
    .Z(_1856_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4331_ (.I(_1856_),
    .ZN(_1857_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4332_ (.A1(_1580_),
    .A2(_1857_),
    .ZN(_1858_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4333_ (.A1(_1761_),
    .A2(_1855_),
    .B(_1858_),
    .ZN(_1859_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4334_ (.I(\soc.spi_video_ram_1.write_fifo.fifo_mem[1][13] ),
    .ZN(_1860_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4335_ (.A1(_1593_),
    .A2(_1860_),
    .B(_1590_),
    .ZN(_1861_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4336_ (.A1(_1756_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[0][13] ),
    .B(_1861_),
    .ZN(_1862_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4337_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[2][13] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[3][13] ),
    .S(_1582_),
    .Z(_1863_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4338_ (.A1(_1710_),
    .A2(_1863_),
    .B(_1579_),
    .ZN(_1864_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4339_ (.A1(_1862_),
    .A2(_1864_),
    .ZN(_1865_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4340_ (.I(\soc.spi_video_ram_1.write_fifo.fifo_mem[5][13] ),
    .ZN(_1866_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4341_ (.A1(_1593_),
    .A2(_1866_),
    .ZN(_1867_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4342_ (.A1(_1756_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[4][13] ),
    .B(_1867_),
    .ZN(_1868_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4343_ (.I(\soc.spi_video_ram_1.write_fifo.fifo_mem[7][13] ),
    .ZN(_1869_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4344_ (.A1(_1755_),
    .A2(_1869_),
    .ZN(_1870_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4345_ (.A1(_1600_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[6][13] ),
    .B(_1870_),
    .C(_1590_),
    .ZN(_1871_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4346_ (.A1(_1591_),
    .A2(_1868_),
    .B(_1871_),
    .C(_1579_),
    .ZN(_1872_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4347_ (.A1(_0703_),
    .A2(_1865_),
    .A3(_1872_),
    .ZN(_1873_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4348_ (.A1(_0686_),
    .A2(_1859_),
    .B1(_1873_),
    .B2(_1850_),
    .ZN(_1874_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4349_ (.A1(_0729_),
    .A2(_1181_),
    .B(_1874_),
    .ZN(_1875_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4350_ (.A1(\soc.spi_video_ram_1.output_buffer[10] ),
    .A2(_1612_),
    .ZN(_1876_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4351_ (.A1(_1811_),
    .A2(_1875_),
    .B(_1876_),
    .ZN(_0070_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4352_ (.I(_1331_),
    .ZN(_1877_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4353_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[0][24] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[1][24] ),
    .I2(\soc.spi_video_ram_1.write_fifo.fifo_mem[2][24] ),
    .I3(\soc.spi_video_ram_1.write_fifo.fifo_mem[3][24] ),
    .S0(_1755_),
    .S1(_1590_),
    .Z(_1878_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4354_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[4][24] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[5][24] ),
    .I2(\soc.spi_video_ram_1.write_fifo.fifo_mem[6][24] ),
    .I3(\soc.spi_video_ram_1.write_fifo.fifo_mem[7][24] ),
    .S0(_1582_),
    .S1(_0001_),
    .Z(_1879_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4355_ (.I(_1879_),
    .ZN(_1880_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4356_ (.A1(_1580_),
    .A2(_1880_),
    .ZN(_1881_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4357_ (.A1(_1761_),
    .A2(_1878_),
    .B(_1881_),
    .ZN(_1882_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4358_ (.I(\soc.spi_video_ram_1.write_fifo.fifo_mem[1][14] ),
    .ZN(_1883_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4359_ (.A1(_1593_),
    .A2(_1883_),
    .B(_1590_),
    .ZN(_1884_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4360_ (.A1(_1756_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[0][14] ),
    .B(_1884_),
    .ZN(_1885_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4361_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[2][14] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[3][14] ),
    .S(_1582_),
    .Z(_1886_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4362_ (.A1(_1710_),
    .A2(_1886_),
    .B(_1579_),
    .ZN(_1887_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4363_ (.A1(_1885_),
    .A2(_1887_),
    .ZN(_1888_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4364_ (.I(\soc.spi_video_ram_1.write_fifo.fifo_mem[5][14] ),
    .ZN(_1889_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4365_ (.A1(_1593_),
    .A2(_1889_),
    .ZN(_1890_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4366_ (.A1(_1600_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[4][14] ),
    .B(_1890_),
    .ZN(_1891_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4367_ (.I(\soc.spi_video_ram_1.write_fifo.fifo_mem[7][14] ),
    .ZN(_1892_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4368_ (.A1(_1755_),
    .A2(_1892_),
    .ZN(_1893_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4369_ (.A1(_1584_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[6][14] ),
    .B(_1893_),
    .C(_1590_),
    .ZN(_1894_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4370_ (.A1(_1710_),
    .A2(_1891_),
    .B(_1894_),
    .C(_1579_),
    .ZN(_1895_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4371_ (.A1(_0703_),
    .A2(_1888_),
    .A3(_1895_),
    .ZN(_1896_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4372_ (.A1(_0686_),
    .A2(_1882_),
    .B1(_1896_),
    .B2(_1850_),
    .ZN(_1897_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4373_ (.A1(_0729_),
    .A2(_1877_),
    .B(_1897_),
    .ZN(_1898_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4374_ (.A1(\soc.spi_video_ram_1.output_buffer[9] ),
    .A2(_1612_),
    .ZN(_1899_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4375_ (.A1(_1811_),
    .A2(_1898_),
    .B(_1899_),
    .ZN(_0071_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4376_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[0][15] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[1][15] ),
    .I2(\soc.spi_video_ram_1.write_fifo.fifo_mem[2][15] ),
    .I3(\soc.spi_video_ram_1.write_fifo.fifo_mem[3][15] ),
    .S0(_1724_),
    .S1(_1587_),
    .Z(_1900_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4377_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[4][15] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[5][15] ),
    .I2(\soc.spi_video_ram_1.write_fifo.fifo_mem[6][15] ),
    .I3(\soc.spi_video_ram_1.write_fifo.fifo_mem[7][15] ),
    .S0(_1583_),
    .S1(_1586_),
    .Z(_1901_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4378_ (.I(_1901_),
    .ZN(_1902_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4379_ (.A1(_1761_),
    .A2(_1902_),
    .ZN(_1903_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4380_ (.A1(_1702_),
    .A2(_1900_),
    .B(_1903_),
    .ZN(_1904_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4381_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[0][23] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[1][23] ),
    .I2(\soc.spi_video_ram_1.write_fifo.fifo_mem[2][23] ),
    .I3(\soc.spi_video_ram_1.write_fifo.fifo_mem[3][23] ),
    .S0(_1755_),
    .S1(_1587_),
    .Z(_1905_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4382_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[4][23] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[5][23] ),
    .I2(\soc.spi_video_ram_1.write_fifo.fifo_mem[6][23] ),
    .I3(\soc.spi_video_ram_1.write_fifo.fifo_mem[7][23] ),
    .S0(_1582_),
    .S1(_0001_),
    .Z(_1906_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4383_ (.I(_1906_),
    .ZN(_1907_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4384_ (.A1(_1580_),
    .A2(_1907_),
    .ZN(_1908_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4385_ (.A1(_1761_),
    .A2(_1905_),
    .B(_1908_),
    .ZN(_1909_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4386_ (.A1(\soc.video_generator_1.v_count[2] ),
    .A2(_1129_),
    .B(_0729_),
    .ZN(_1910_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _4387_ (.A1(_1821_),
    .A2(_1904_),
    .B1(_1909_),
    .B2(_1850_),
    .C(_1910_),
    .ZN(_1911_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4388_ (.A1(\soc.spi_video_ram_1.output_buffer[8] ),
    .A2(_1612_),
    .B1(_1825_),
    .B2(_1911_),
    .ZN(_1912_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4389_ (.I(_1912_),
    .ZN(_0072_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4390_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[0][22] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[1][22] ),
    .S(_1584_),
    .Z(_1913_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4391_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[2][22] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[3][22] ),
    .S(_1584_),
    .Z(_1914_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4392_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[4][22] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[5][22] ),
    .S(_1584_),
    .Z(_1915_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4393_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[6][22] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[7][22] ),
    .S(_1584_),
    .Z(_1916_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4394_ (.I0(_1913_),
    .I1(_1914_),
    .I2(_1915_),
    .I3(_1916_),
    .S0(_1591_),
    .S1(_1761_),
    .Z(_1917_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4395_ (.A1(_1144_),
    .A2(_1695_),
    .ZN(_1918_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4396_ (.A1(_1609_),
    .A2(_1917_),
    .B(_1918_),
    .ZN(_1919_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4397_ (.A1(\soc.spi_video_ram_1.output_buffer[7] ),
    .A2(_1611_),
    .ZN(_1920_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4398_ (.A1(_1686_),
    .A2(_1919_),
    .B(_1920_),
    .ZN(_0073_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4399_ (.I(_1695_),
    .ZN(_1921_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4400_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[0][21] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[1][21] ),
    .S(_1724_),
    .Z(_1922_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4401_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[2][21] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[3][21] ),
    .S(_1724_),
    .Z(_1923_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4402_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[4][21] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[5][21] ),
    .S(_1724_),
    .Z(_1924_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4403_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[6][21] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[7][21] ),
    .S(_1724_),
    .Z(_1925_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4404_ (.I0(_1922_),
    .I1(_1923_),
    .I2(_1924_),
    .I3(_1925_),
    .S0(_1710_),
    .S1(_1580_),
    .Z(_1926_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4405_ (.A1(_1140_),
    .A2(_1921_),
    .B1(_1926_),
    .B2(_1609_),
    .ZN(_1927_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4406_ (.A1(\soc.spi_video_ram_1.output_buffer[6] ),
    .A2(_1611_),
    .ZN(_1928_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4407_ (.A1(_1686_),
    .A2(_1927_),
    .B(_1928_),
    .ZN(_0074_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4408_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[0][20] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[1][20] ),
    .I2(\soc.spi_video_ram_1.write_fifo.fifo_mem[2][20] ),
    .I3(\soc.spi_video_ram_1.write_fifo.fifo_mem[3][20] ),
    .S0(_1594_),
    .S1(_1588_),
    .Z(_1929_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4409_ (.I(\soc.spi_video_ram_1.write_fifo.fifo_mem[5][20] ),
    .ZN(_1930_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4410_ (.A1(_1585_),
    .A2(_1930_),
    .ZN(_1931_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4411_ (.A1(_1601_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[4][20] ),
    .B(_1931_),
    .ZN(_1932_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4412_ (.I(\soc.spi_video_ram_1.write_fifo.fifo_mem[7][20] ),
    .ZN(_1933_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4413_ (.A1(_1756_),
    .A2(_1933_),
    .ZN(_1934_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4414_ (.A1(_1596_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[6][20] ),
    .B(_1934_),
    .C(_1591_),
    .ZN(_1935_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4415_ (.A1(_1592_),
    .A2(_1932_),
    .B(_1935_),
    .C(_1702_),
    .ZN(_1936_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4416_ (.A1(_1581_),
    .A2(_1929_),
    .B(_1936_),
    .C(_1609_),
    .ZN(_1937_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4417_ (.A1(\soc.spi_video_ram_1.output_buffer[5] ),
    .A2(_1611_),
    .ZN(_1938_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4418_ (.A1(_1578_),
    .A2(_1937_),
    .B(_1938_),
    .ZN(_0075_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4419_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[0][19] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[1][19] ),
    .I2(\soc.spi_video_ram_1.write_fifo.fifo_mem[2][19] ),
    .I3(\soc.spi_video_ram_1.write_fifo.fifo_mem[3][19] ),
    .S0(_1594_),
    .S1(_1588_),
    .Z(_1939_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4420_ (.I(\soc.spi_video_ram_1.write_fifo.fifo_mem[5][19] ),
    .ZN(_1940_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4421_ (.A1(_1585_),
    .A2(_1940_),
    .ZN(_1941_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4422_ (.A1(_1601_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[4][19] ),
    .B(_1941_),
    .ZN(_1942_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4423_ (.I(\soc.spi_video_ram_1.write_fifo.fifo_mem[7][19] ),
    .ZN(_1943_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4424_ (.A1(_1756_),
    .A2(_1943_),
    .ZN(_1944_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4425_ (.A1(_1596_),
    .A2(\soc.spi_video_ram_1.write_fifo.fifo_mem[6][19] ),
    .B(_1944_),
    .C(_1591_),
    .ZN(_1945_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4426_ (.A1(_1592_),
    .A2(_1942_),
    .B(_1945_),
    .C(_1702_),
    .ZN(_1946_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4427_ (.A1(_1581_),
    .A2(_1939_),
    .B(_1946_),
    .C(_1609_),
    .ZN(_1947_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4428_ (.A1(\soc.spi_video_ram_1.output_buffer[4] ),
    .A2(_1611_),
    .ZN(_1948_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4429_ (.A1(_1578_),
    .A2(_1947_),
    .B(_1948_),
    .ZN(_0076_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4430_ (.I(\soc.spi_video_ram_1.fifo_read_request ),
    .ZN(_1949_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4431_ (.A1(_1949_),
    .A2(_0702_),
    .ZN(_1950_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4432_ (.A1(\soc.spi_video_ram_1.write_fifo.read_pointer[0] ),
    .A2(_1950_),
    .ZN(_1951_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _4433_ (.A1(_0697_),
    .A2(_1949_),
    .A3(_0702_),
    .ZN(_1952_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _4434_ (.A1(_1461_),
    .A2(_1951_),
    .A3(_1952_),
    .ZN(_0077_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4435_ (.A1(\soc.spi_video_ram_1.write_fifo.read_pointer[1] ),
    .A2(_1952_),
    .ZN(_1953_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4436_ (.A1(\soc.spi_video_ram_1.write_fifo.read_pointer[1] ),
    .A2(_1952_),
    .Z(_1954_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _4437_ (.A1(_1461_),
    .A2(_1953_),
    .A3(_1954_),
    .ZN(_0078_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4438_ (.I(_0675_),
    .Z(_1955_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4439_ (.A1(\soc.spi_video_ram_1.write_fifo.read_pointer[2] ),
    .A2(_1954_),
    .Z(_1956_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4440_ (.A1(_1955_),
    .A2(_1956_),
    .Z(_1957_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4441_ (.I(_1957_),
    .Z(_0079_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4442_ (.A1(_0708_),
    .A2(_0705_),
    .B1(_0732_),
    .B2(\soc.spi_video_ram_1.current_state[4] ),
    .ZN(_1958_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _4443_ (.A1(_0688_),
    .A2(_0726_),
    .A3(_0735_),
    .A4(_1958_),
    .ZN(_1959_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4444_ (.A1(_0709_),
    .A2(_1959_),
    .B(_0674_),
    .ZN(_1960_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4445_ (.I(_1960_),
    .Z(_1961_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4446_ (.A1(\soc.spi_video_ram_1.state_counter[0] ),
    .A2(_1961_),
    .ZN(_0080_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4447_ (.A1(\soc.spi_video_ram_1.state_counter[1] ),
    .A2(\soc.spi_video_ram_1.state_counter[0] ),
    .ZN(_1962_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4448_ (.A1(_1961_),
    .A2(_1962_),
    .ZN(_0081_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _4449_ (.A1(\soc.spi_video_ram_1.state_counter[1] ),
    .A2(\soc.spi_video_ram_1.state_counter[0] ),
    .A3(\soc.spi_video_ram_1.state_counter[2] ),
    .Z(_1963_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4450_ (.A1(\soc.spi_video_ram_1.state_counter[1] ),
    .A2(\soc.spi_video_ram_1.state_counter[0] ),
    .B(\soc.spi_video_ram_1.state_counter[2] ),
    .ZN(_1964_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _4451_ (.A1(_1961_),
    .A2(_1963_),
    .A3(_1964_),
    .ZN(_0082_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4452_ (.A1(\soc.spi_video_ram_1.state_counter[3] ),
    .A2(_1963_),
    .Z(_1965_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4453_ (.A1(\soc.spi_video_ram_1.state_counter[3] ),
    .A2(_1963_),
    .ZN(_1966_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _4454_ (.A1(_1961_),
    .A2(_1965_),
    .A3(_1966_),
    .ZN(_0083_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4455_ (.A1(\soc.spi_video_ram_1.state_counter[4] ),
    .A2(_1965_),
    .Z(_1967_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4456_ (.A1(\soc.spi_video_ram_1.state_counter[4] ),
    .A2(_1965_),
    .ZN(_1968_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _4457_ (.A1(_1961_),
    .A2(_1967_),
    .A3(_1968_),
    .ZN(_0084_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4458_ (.A1(\soc.spi_video_ram_1.state_counter[5] ),
    .A2(_1967_),
    .Z(_1969_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4459_ (.A1(\soc.spi_video_ram_1.state_counter[5] ),
    .A2(_1967_),
    .ZN(_1970_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _4460_ (.A1(_1961_),
    .A2(_1969_),
    .A3(_1970_),
    .ZN(_0085_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4461_ (.A1(\soc.spi_video_ram_1.state_counter[6] ),
    .A2(_1969_),
    .Z(_1971_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4462_ (.A1(\soc.spi_video_ram_1.state_counter[6] ),
    .A2(_1969_),
    .ZN(_1972_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _4463_ (.A1(_1961_),
    .A2(_1971_),
    .A3(_1972_),
    .ZN(_0086_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4464_ (.A1(\soc.spi_video_ram_1.state_counter[7] ),
    .A2(_1971_),
    .Z(_1973_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4465_ (.A1(\soc.spi_video_ram_1.state_counter[7] ),
    .A2(_1971_),
    .ZN(_1974_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _4466_ (.A1(_1961_),
    .A2(_1973_),
    .A3(_1974_),
    .ZN(_0087_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4467_ (.A1(\soc.spi_video_ram_1.state_counter[8] ),
    .A2(_1973_),
    .Z(_1975_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4468_ (.A1(\soc.spi_video_ram_1.state_counter[8] ),
    .A2(_1973_),
    .ZN(_1976_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _4469_ (.A1(_1960_),
    .A2(_1975_),
    .A3(_1976_),
    .ZN(_0088_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4470_ (.A1(\soc.spi_video_ram_1.state_counter[9] ),
    .A2(_1975_),
    .ZN(_1977_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4471_ (.A1(_1961_),
    .A2(_1977_),
    .ZN(_0089_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4472_ (.A1(\soc.spi_video_ram_1.state_counter[9] ),
    .A2(_1975_),
    .ZN(_1978_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4473_ (.A1(\soc.spi_video_ram_1.state_counter[10] ),
    .A2(_1978_),
    .Z(_1979_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4474_ (.A1(_1961_),
    .A2(_1979_),
    .ZN(_0090_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4475_ (.A1(\soc.video_generator_1.v_count[0] ),
    .A2(_1458_),
    .Z(_1980_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _4476_ (.A1(_1125_),
    .A2(\soc.video_generator_1.v_count[8] ),
    .A3(\soc.video_generator_1.v_count[7] ),
    .A4(_1126_),
    .ZN(_1981_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _4477_ (.A1(_1162_),
    .A2(\soc.video_generator_1.v_count[1] ),
    .A3(_1139_),
    .ZN(_1982_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _4478_ (.A1(\soc.video_generator_1.v_count[2] ),
    .A2(_1981_),
    .A3(_1982_),
    .ZN(_1983_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_4 _4479_ (.A1(_1127_),
    .A2(_1167_),
    .A3(_1983_),
    .B(_0675_),
    .ZN(_1984_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4480_ (.A1(\soc.video_generator_1.v_count[0] ),
    .A2(_1458_),
    .ZN(_1985_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _4481_ (.A1(_1980_),
    .A2(_1984_),
    .A3(_1985_),
    .ZN(_0091_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4482_ (.A1(\soc.video_generator_1.v_count[1] ),
    .A2(_1980_),
    .ZN(_1986_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4483_ (.A1(\soc.video_generator_1.v_count[1] ),
    .A2(_1980_),
    .Z(_1987_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _4484_ (.A1(_1984_),
    .A2(_1986_),
    .A3(_1987_),
    .ZN(_0092_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4485_ (.A1(\soc.video_generator_1.v_count[2] ),
    .A2(_1987_),
    .ZN(_1988_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4486_ (.A1(\soc.video_generator_1.v_count[2] ),
    .A2(_1987_),
    .Z(_1989_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _4487_ (.A1(_1984_),
    .A2(_1988_),
    .A3(_1989_),
    .ZN(_0093_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4488_ (.A1(\soc.video_generator_1.v_count[3] ),
    .A2(_1989_),
    .ZN(_1990_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4489_ (.A1(\soc.video_generator_1.v_count[3] ),
    .A2(_1989_),
    .Z(_1991_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _4490_ (.A1(_1984_),
    .A2(_1990_),
    .A3(_1991_),
    .ZN(_0094_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4491_ (.A1(_1167_),
    .A2(_1991_),
    .ZN(_1992_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4492_ (.A1(_1167_),
    .A2(_1991_),
    .Z(_1993_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _4493_ (.A1(_1984_),
    .A2(_1992_),
    .A3(_1993_),
    .ZN(_0095_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4494_ (.A1(_1127_),
    .A2(_1993_),
    .ZN(_1994_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4495_ (.A1(_1127_),
    .A2(_1993_),
    .Z(_1995_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _4496_ (.A1(_1984_),
    .A2(_1994_),
    .A3(_1995_),
    .ZN(_0096_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4497_ (.A1(_1126_),
    .A2(_1995_),
    .ZN(_1996_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _4498_ (.A1(_1126_),
    .A2(_1995_),
    .B(_1996_),
    .C(_1984_),
    .ZN(_0097_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4499_ (.A1(_1126_),
    .A2(_1995_),
    .B(\soc.video_generator_1.v_count[7] ),
    .ZN(_1997_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4500_ (.A1(_1167_),
    .A2(_1991_),
    .ZN(_1998_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4501_ (.A1(_1168_),
    .A2(_1998_),
    .ZN(_1999_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _4502_ (.A1(_1984_),
    .A2(_1997_),
    .A3(_1999_),
    .ZN(_0098_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4503_ (.A1(\soc.video_generator_1.v_count[8] ),
    .A2(_1999_),
    .ZN(_2000_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4504_ (.A1(_1128_),
    .A2(_1998_),
    .ZN(_2001_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _4505_ (.A1(_1984_),
    .A2(_2000_),
    .A3(_2001_),
    .ZN(_0099_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4506_ (.A1(_1142_),
    .A2(_2001_),
    .ZN(_2002_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _4507_ (.A1(_1142_),
    .A2(_2001_),
    .B(_2002_),
    .C(_1984_),
    .ZN(_0100_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4508_ (.I(_0748_),
    .Z(_2003_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4509_ (.A1(\soc.spi_video_ram_1.fifo_in_data[0] ),
    .A2(_2003_),
    .ZN(_2004_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4510_ (.A1(_0009_),
    .A2(_0878_),
    .B(_2004_),
    .ZN(_0101_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4511_ (.A1(\soc.spi_video_ram_1.fifo_in_data[1] ),
    .A2(_2003_),
    .ZN(_2005_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4512_ (.A1(_0009_),
    .A2(_0902_),
    .B(_2005_),
    .ZN(_0102_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4513_ (.A1(\soc.spi_video_ram_1.fifo_in_data[2] ),
    .A2(_2003_),
    .ZN(_2006_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4514_ (.A1(_0009_),
    .A2(_0920_),
    .B(_2006_),
    .ZN(_0103_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4515_ (.I(_0748_),
    .Z(_2007_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4516_ (.A1(\soc.spi_video_ram_1.fifo_in_data[3] ),
    .A2(_2007_),
    .ZN(_2008_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4517_ (.A1(_0009_),
    .A2(_0942_),
    .B(_2008_),
    .ZN(_0104_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4518_ (.A1(\soc.spi_video_ram_1.fifo_in_data[4] ),
    .A2(_2007_),
    .ZN(_2009_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4519_ (.A1(_0009_),
    .A2(_0958_),
    .B(_2009_),
    .ZN(_0105_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4520_ (.A1(\soc.spi_video_ram_1.fifo_in_data[5] ),
    .A2(_2007_),
    .ZN(_2010_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4521_ (.A1(_0009_),
    .A2(_0970_),
    .B(_2010_),
    .ZN(_0106_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4522_ (.A1(\soc.spi_video_ram_1.fifo_in_data[6] ),
    .A2(_2007_),
    .ZN(_2011_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4523_ (.A1(_0009_),
    .A2(_0989_),
    .B(_2011_),
    .ZN(_0107_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4524_ (.A1(\soc.spi_video_ram_1.fifo_in_data[7] ),
    .A2(_2007_),
    .ZN(_2012_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4525_ (.A1(_0009_),
    .A2(_1002_),
    .B(_2012_),
    .ZN(_0108_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4526_ (.A1(\soc.spi_video_ram_1.fifo_in_data[8] ),
    .A2(_2007_),
    .ZN(_2013_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4527_ (.A1(_0009_),
    .A2(_1024_),
    .B(_2013_),
    .ZN(_0109_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4528_ (.A1(\soc.spi_video_ram_1.fifo_in_data[9] ),
    .A2(_2007_),
    .ZN(_2014_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4529_ (.A1(_2003_),
    .A2(_1039_),
    .B(_2014_),
    .ZN(_0110_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4530_ (.A1(\soc.spi_video_ram_1.fifo_in_data[10] ),
    .A2(_2007_),
    .ZN(_2015_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4531_ (.A1(_2003_),
    .A2(_1058_),
    .B(_2015_),
    .ZN(_0111_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4532_ (.A1(\soc.spi_video_ram_1.fifo_in_data[11] ),
    .A2(_2007_),
    .ZN(_2016_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4533_ (.A1(_2003_),
    .A2(_1069_),
    .B(_2016_),
    .ZN(_0112_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4534_ (.A1(\soc.spi_video_ram_1.fifo_in_data[12] ),
    .A2(_2007_),
    .ZN(_2017_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4535_ (.A1(_2003_),
    .A2(_1092_),
    .B(_2017_),
    .ZN(_0113_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 _4536_ (.I(_0748_),
    .Z(_2018_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4537_ (.A1(\soc.spi_video_ram_1.fifo_in_data[13] ),
    .A2(_2018_),
    .ZN(_2019_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4538_ (.A1(_2003_),
    .A2(_1108_),
    .B(_2019_),
    .ZN(_0114_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4539_ (.A1(\soc.spi_video_ram_1.fifo_in_data[14] ),
    .A2(_2018_),
    .ZN(_2020_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4540_ (.A1(_2003_),
    .A2(_1123_),
    .B(_2020_),
    .ZN(_0115_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4541_ (.A1(\soc.spi_video_ram_1.fifo_in_data[15] ),
    .A2(_2018_),
    .ZN(_2021_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4542_ (.A1(_2003_),
    .A2(_1669_),
    .B(_2021_),
    .ZN(_0116_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _4543_ (.A1(\soc.spi_video_ram_1.write_fifo.write_pointer[2] ),
    .A2(_0694_),
    .A3(_0698_),
    .ZN(_2022_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 _4544_ (.I(_2022_),
    .Z(_2023_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4545_ (.I0(\soc.spi_video_ram_1.fifo_in_data[0] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[7][0] ),
    .S(_2023_),
    .Z(_2024_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4546_ (.I(_2024_),
    .Z(_0117_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4547_ (.I(_2022_),
    .Z(_2025_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4548_ (.I(_2022_),
    .Z(_2026_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4549_ (.A1(\soc.spi_video_ram_1.fifo_in_data[1] ),
    .A2(_2026_),
    .ZN(_2027_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4550_ (.A1(_1708_),
    .A2(_2025_),
    .B(_2027_),
    .ZN(_0118_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4551_ (.I0(\soc.spi_video_ram_1.fifo_in_data[2] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[7][2] ),
    .S(_2023_),
    .Z(_2028_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4552_ (.I(_2028_),
    .Z(_0119_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4553_ (.I0(\soc.spi_video_ram_1.fifo_in_data[3] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[7][3] ),
    .S(_2023_),
    .Z(_2029_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4554_ (.I(_2029_),
    .Z(_0120_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4555_ (.I0(\soc.spi_video_ram_1.fifo_in_data[4] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[7][4] ),
    .S(_2023_),
    .Z(_2030_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4556_ (.I(_2030_),
    .Z(_0121_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4557_ (.A1(\soc.spi_video_ram_1.fifo_in_data[5] ),
    .A2(_2026_),
    .ZN(_2031_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4558_ (.A1(_1743_),
    .A2(_2025_),
    .B(_2031_),
    .ZN(_0122_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4559_ (.A1(\soc.spi_video_ram_1.fifo_in_data[6] ),
    .A2(_2026_),
    .ZN(_2032_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4560_ (.A1(_1757_),
    .A2(_2025_),
    .B(_2032_),
    .ZN(_0123_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4561_ (.A1(\soc.spi_video_ram_1.fifo_in_data[7] ),
    .A2(_2026_),
    .ZN(_2033_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4562_ (.A1(_1770_),
    .A2(_2025_),
    .B(_2033_),
    .ZN(_0124_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4563_ (.A1(\soc.spi_video_ram_1.fifo_in_data[8] ),
    .A2(_2026_),
    .ZN(_2034_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4564_ (.A1(_1790_),
    .A2(_2025_),
    .B(_2034_),
    .ZN(_0125_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4565_ (.I0(\soc.spi_video_ram_1.fifo_in_data[9] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[7][9] ),
    .S(_2023_),
    .Z(_2035_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4566_ (.I(_2035_),
    .Z(_0126_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4567_ (.I0(\soc.spi_video_ram_1.fifo_in_data[10] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[7][10] ),
    .S(_2023_),
    .Z(_2036_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4568_ (.I(_2036_),
    .Z(_0127_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _4569_ (.I(_2022_),
    .Z(_2037_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4570_ (.I0(\soc.spi_video_ram_1.fifo_in_data[11] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[7][11] ),
    .S(_2037_),
    .Z(_2038_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4571_ (.I(_2038_),
    .Z(_0128_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4572_ (.I0(\soc.spi_video_ram_1.fifo_in_data[12] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[7][12] ),
    .S(_2037_),
    .Z(_2039_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4573_ (.I(_2039_),
    .Z(_0129_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4574_ (.A1(\soc.spi_video_ram_1.fifo_in_data[13] ),
    .A2(_2026_),
    .ZN(_2040_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4575_ (.A1(_1869_),
    .A2(_2025_),
    .B(_2040_),
    .ZN(_0130_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4576_ (.A1(\soc.spi_video_ram_1.fifo_in_data[14] ),
    .A2(_2026_),
    .ZN(_2041_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4577_ (.A1(_1892_),
    .A2(_2025_),
    .B(_2041_),
    .ZN(_0131_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4578_ (.I0(\soc.spi_video_ram_1.fifo_in_data[15] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[7][15] ),
    .S(_2037_),
    .Z(_2042_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4579_ (.I(_2042_),
    .Z(_0132_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4580_ (.A1(\soc.spi_video_ram_1.fifo_in_address[0] ),
    .A2(_2026_),
    .ZN(_2043_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4581_ (.A1(_1602_),
    .A2(_2025_),
    .B(_2043_),
    .ZN(_0133_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4582_ (.A1(\soc.spi_video_ram_1.fifo_in_address[1] ),
    .A2(_2023_),
    .ZN(_2044_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4583_ (.A1(_1628_),
    .A2(_2025_),
    .B(_2044_),
    .ZN(_0134_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4584_ (.A1(\soc.spi_video_ram_1.fifo_in_address[2] ),
    .A2(_2023_),
    .ZN(_2045_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4585_ (.A1(_1618_),
    .A2(_2025_),
    .B(_2045_),
    .ZN(_0135_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4586_ (.A1(\soc.spi_video_ram_1.fifo_in_address[3] ),
    .A2(_2023_),
    .ZN(_2046_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4587_ (.A1(_1943_),
    .A2(_2026_),
    .B(_2046_),
    .ZN(_0136_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4588_ (.A1(\soc.spi_video_ram_1.fifo_in_address[4] ),
    .A2(_2023_),
    .ZN(_2047_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4589_ (.A1(_1933_),
    .A2(_2026_),
    .B(_2047_),
    .ZN(_0137_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4590_ (.I0(\soc.spi_video_ram_1.fifo_in_address[5] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[7][21] ),
    .S(_2037_),
    .Z(_2048_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4591_ (.I(_2048_),
    .Z(_0138_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4592_ (.I0(\soc.spi_video_ram_1.fifo_in_address[6] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[7][22] ),
    .S(_2037_),
    .Z(_2049_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4593_ (.I(_2049_),
    .Z(_0139_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4594_ (.I0(\soc.spi_video_ram_1.fifo_in_address[7] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[7][23] ),
    .S(_2037_),
    .Z(_2050_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4595_ (.I(_2050_),
    .Z(_0140_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4596_ (.I0(\soc.spi_video_ram_1.fifo_in_address[8] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[7][24] ),
    .S(_2037_),
    .Z(_2051_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4597_ (.I(_2051_),
    .Z(_0141_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4598_ (.I0(\soc.spi_video_ram_1.fifo_in_address[9] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[7][25] ),
    .S(_2037_),
    .Z(_2052_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4599_ (.I(_2052_),
    .Z(_0142_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4600_ (.I0(\soc.spi_video_ram_1.fifo_in_address[10] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[7][26] ),
    .S(_2037_),
    .Z(_2053_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4601_ (.I(_2053_),
    .Z(_0143_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4602_ (.I0(\soc.spi_video_ram_1.fifo_in_address[11] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[7][27] ),
    .S(_2037_),
    .Z(_2054_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4603_ (.I(_2054_),
    .Z(_0144_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4604_ (.I0(\soc.spi_video_ram_1.fifo_in_address[12] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[7][28] ),
    .S(_2022_),
    .Z(_2055_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4605_ (.I(_2055_),
    .Z(_0145_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _4606_ (.A1(_0700_),
    .A2(_0694_),
    .A3(_0698_),
    .ZN(_2056_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _4607_ (.I(_2056_),
    .Z(_2057_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _4608_ (.I(_2057_),
    .Z(_2058_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4609_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[4][0] ),
    .I1(\soc.spi_video_ram_1.fifo_in_data[0] ),
    .S(_2058_),
    .Z(_2059_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4610_ (.I(_2059_),
    .Z(_0146_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4611_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[4][1] ),
    .I1(\soc.spi_video_ram_1.fifo_in_data[1] ),
    .S(_2058_),
    .Z(_2060_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4612_ (.I(_2060_),
    .Z(_0147_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4613_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[4][2] ),
    .I1(\soc.spi_video_ram_1.fifo_in_data[2] ),
    .S(_2058_),
    .Z(_2061_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4614_ (.I(_2061_),
    .Z(_0148_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4615_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[4][3] ),
    .I1(\soc.spi_video_ram_1.fifo_in_data[3] ),
    .S(_2058_),
    .Z(_2062_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4616_ (.I(_2062_),
    .Z(_0149_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4617_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[4][4] ),
    .I1(\soc.spi_video_ram_1.fifo_in_data[4] ),
    .S(_2058_),
    .Z(_2063_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4618_ (.I(_2063_),
    .Z(_0150_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4619_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[4][5] ),
    .I1(\soc.spi_video_ram_1.fifo_in_data[5] ),
    .S(_2058_),
    .Z(_2064_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4620_ (.I(_2064_),
    .Z(_0151_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4621_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[4][6] ),
    .I1(\soc.spi_video_ram_1.fifo_in_data[6] ),
    .S(_2058_),
    .Z(_2065_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4622_ (.I(_2065_),
    .Z(_0152_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4623_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[4][7] ),
    .I1(\soc.spi_video_ram_1.fifo_in_data[7] ),
    .S(_2058_),
    .Z(_2066_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4624_ (.I(_2066_),
    .Z(_0153_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4625_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[4][8] ),
    .I1(\soc.spi_video_ram_1.fifo_in_data[8] ),
    .S(_2058_),
    .Z(_2067_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4626_ (.I(_2067_),
    .Z(_0154_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4627_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[4][9] ),
    .I1(\soc.spi_video_ram_1.fifo_in_data[9] ),
    .S(_2058_),
    .Z(_2068_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4628_ (.I(_2068_),
    .Z(_0155_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _4629_ (.I(_2056_),
    .Z(_2069_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4630_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[4][10] ),
    .I1(\soc.spi_video_ram_1.fifo_in_data[10] ),
    .S(_2069_),
    .Z(_2070_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4631_ (.I(_2070_),
    .Z(_0156_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4632_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[4][11] ),
    .I1(\soc.spi_video_ram_1.fifo_in_data[11] ),
    .S(_2069_),
    .Z(_2071_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4633_ (.I(_2071_),
    .Z(_0157_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4634_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[4][12] ),
    .I1(\soc.spi_video_ram_1.fifo_in_data[12] ),
    .S(_2069_),
    .Z(_2072_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4635_ (.I(_2072_),
    .Z(_0158_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4636_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[4][13] ),
    .I1(\soc.spi_video_ram_1.fifo_in_data[13] ),
    .S(_2069_),
    .Z(_2073_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4637_ (.I(_2073_),
    .Z(_0159_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4638_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[4][14] ),
    .I1(\soc.spi_video_ram_1.fifo_in_data[14] ),
    .S(_2069_),
    .Z(_2074_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4639_ (.I(_2074_),
    .Z(_0160_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4640_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[4][15] ),
    .I1(\soc.spi_video_ram_1.fifo_in_data[15] ),
    .S(_2069_),
    .Z(_2075_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4641_ (.I(_2075_),
    .Z(_0161_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4642_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[4][16] ),
    .I1(\soc.spi_video_ram_1.fifo_in_address[0] ),
    .S(_2069_),
    .Z(_2076_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4643_ (.I(_2076_),
    .Z(_0162_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4644_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[4][17] ),
    .I1(\soc.spi_video_ram_1.fifo_in_address[1] ),
    .S(_2069_),
    .Z(_2077_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4645_ (.I(_2077_),
    .Z(_0163_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4646_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[4][18] ),
    .I1(\soc.spi_video_ram_1.fifo_in_address[2] ),
    .S(_2069_),
    .Z(_2078_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4647_ (.I(_2078_),
    .Z(_0164_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4648_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[4][19] ),
    .I1(\soc.spi_video_ram_1.fifo_in_address[3] ),
    .S(_2069_),
    .Z(_2079_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4649_ (.I(_2079_),
    .Z(_0165_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4650_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[4][20] ),
    .I1(\soc.spi_video_ram_1.fifo_in_address[4] ),
    .S(_2057_),
    .Z(_2080_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4651_ (.I(_2080_),
    .Z(_0166_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4652_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[4][21] ),
    .I1(\soc.spi_video_ram_1.fifo_in_address[5] ),
    .S(_2057_),
    .Z(_2081_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4653_ (.I(_2081_),
    .Z(_0167_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4654_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[4][22] ),
    .I1(\soc.spi_video_ram_1.fifo_in_address[6] ),
    .S(_2057_),
    .Z(_2082_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4655_ (.I(_2082_),
    .Z(_0168_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4656_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[4][23] ),
    .I1(\soc.spi_video_ram_1.fifo_in_address[7] ),
    .S(_2057_),
    .Z(_2083_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4657_ (.I(_2083_),
    .Z(_0169_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4658_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[4][24] ),
    .I1(\soc.spi_video_ram_1.fifo_in_address[8] ),
    .S(_2057_),
    .Z(_2084_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4659_ (.I(_2084_),
    .Z(_0170_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4660_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[4][25] ),
    .I1(\soc.spi_video_ram_1.fifo_in_address[9] ),
    .S(_2057_),
    .Z(_2085_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4661_ (.I(_2085_),
    .Z(_0171_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4662_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[4][26] ),
    .I1(\soc.spi_video_ram_1.fifo_in_address[10] ),
    .S(_2057_),
    .Z(_2086_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4663_ (.I(_2086_),
    .Z(_0172_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4664_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[4][27] ),
    .I1(\soc.spi_video_ram_1.fifo_in_address[11] ),
    .S(_2057_),
    .Z(_2087_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4665_ (.I(_2087_),
    .Z(_0173_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4666_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[4][28] ),
    .I1(\soc.spi_video_ram_1.fifo_in_address[12] ),
    .S(_2057_),
    .Z(_2088_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4667_ (.I(_2088_),
    .Z(_0174_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _4668_ (.I(\soc.rom_encoder_0.write_enable ),
    .ZN(_2089_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4669_ (.A1(_2089_),
    .A2(_0689_),
    .ZN(_2090_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4670_ (.I(_2090_),
    .Z(_0175_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _4671_ (.A1(\soc.spi_video_ram_1.current_state[3] ),
    .A2(_0703_),
    .A3(\soc.spi_video_ram_1.current_state[0] ),
    .A4(\soc.spi_video_ram_1.current_state[2] ),
    .ZN(_2091_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4672_ (.A1(_2091_),
    .A2(_1962_),
    .ZN(_2092_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4673_ (.A1(\soc.spi_video_ram_1.state_counter[0] ),
    .A2(_2091_),
    .B(_2092_),
    .ZN(_2093_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4674_ (.A1(net69),
    .A2(_2093_),
    .ZN(_2094_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4675_ (.A1(\soc.spi_video_ram_1.state_sram_clk_counter[0] ),
    .A2(_2094_),
    .Z(_2095_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _4676_ (.A1(\soc.spi_video_ram_1.current_state[2] ),
    .A2(net68),
    .ZN(_2096_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4677_ (.A1(\soc.spi_video_ram_1.state_sram_clk_counter[0] ),
    .A2(_2094_),
    .B(_2096_),
    .ZN(_2097_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4678_ (.A1(_2095_),
    .A2(_2097_),
    .ZN(_0176_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4679_ (.A1(\soc.spi_video_ram_1.state_sram_clk_counter[1] ),
    .A2(_2095_),
    .Z(_2098_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4680_ (.A1(\soc.spi_video_ram_1.state_sram_clk_counter[1] ),
    .A2(_2095_),
    .B(_2096_),
    .ZN(_2099_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4681_ (.A1(_2098_),
    .A2(_2099_),
    .ZN(_0177_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4682_ (.A1(\soc.spi_video_ram_1.state_sram_clk_counter[2] ),
    .A2(_2098_),
    .Z(_2100_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4683_ (.A1(\soc.spi_video_ram_1.state_sram_clk_counter[2] ),
    .A2(_2098_),
    .B(_2096_),
    .ZN(_2101_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4684_ (.A1(_2100_),
    .A2(_2101_),
    .ZN(_0178_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4685_ (.A1(\soc.spi_video_ram_1.state_sram_clk_counter[3] ),
    .A2(_2100_),
    .Z(_2102_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4686_ (.A1(\soc.spi_video_ram_1.state_sram_clk_counter[3] ),
    .A2(_2100_),
    .B(_2096_),
    .ZN(_2103_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4687_ (.A1(_2102_),
    .A2(_2103_),
    .ZN(_0179_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4688_ (.A1(\soc.spi_video_ram_1.state_sram_clk_counter[4] ),
    .A2(_2102_),
    .Z(_2104_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4689_ (.A1(\soc.spi_video_ram_1.state_sram_clk_counter[4] ),
    .A2(_2102_),
    .B(_2096_),
    .ZN(_2105_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4690_ (.A1(_2104_),
    .A2(_2105_),
    .ZN(_0180_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4691_ (.A1(\soc.spi_video_ram_1.state_sram_clk_counter[5] ),
    .A2(_2104_),
    .Z(_2106_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4692_ (.A1(\soc.spi_video_ram_1.state_sram_clk_counter[5] ),
    .A2(_2104_),
    .B(_2096_),
    .ZN(_2107_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4693_ (.A1(_2106_),
    .A2(_2107_),
    .ZN(_0181_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4694_ (.A1(\soc.spi_video_ram_1.state_sram_clk_counter[6] ),
    .A2(_2106_),
    .Z(_2108_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4695_ (.A1(\soc.spi_video_ram_1.state_sram_clk_counter[6] ),
    .A2(_2106_),
    .B(_2096_),
    .ZN(_2109_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4696_ (.A1(_2108_),
    .A2(_2109_),
    .ZN(_0182_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4697_ (.A1(\soc.spi_video_ram_1.state_sram_clk_counter[7] ),
    .A2(_2108_),
    .B(_2096_),
    .ZN(_2110_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4698_ (.A1(\soc.spi_video_ram_1.state_sram_clk_counter[7] ),
    .A2(_2108_),
    .B(_2110_),
    .ZN(_0183_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4699_ (.A1(\soc.spi_video_ram_1.current_state[2] ),
    .A2(net68),
    .Z(_2111_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4700_ (.A1(\soc.spi_video_ram_1.state_sram_clk_counter[7] ),
    .A2(_2108_),
    .ZN(_2112_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4701_ (.A1(\soc.spi_video_ram_1.state_sram_clk_counter[8] ),
    .A2(_2112_),
    .Z(_2113_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4702_ (.A1(_2111_),
    .A2(_2113_),
    .ZN(_0184_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4703_ (.A1(_2093_),
    .A2(_2111_),
    .ZN(_0185_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _4704_ (.A1(net69),
    .A2(_2093_),
    .A3(_2111_),
    .ZN(_0186_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _4705_ (.A1(net69),
    .A2(_2093_),
    .A3(_2096_),
    .Z(_2114_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4706_ (.I(_2114_),
    .Z(_0187_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4707_ (.A1(\soc.spi_video_ram_1.state_sram_clk_counter[2] ),
    .A2(\soc.spi_video_ram_1.state_sram_clk_counter[1] ),
    .B(\soc.spi_video_ram_1.state_sram_clk_counter[3] ),
    .ZN(_2115_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4708_ (.A1(_0682_),
    .A2(_2115_),
    .ZN(_2116_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _4709_ (.A1(\soc.spi_video_ram_1.state_sram_clk_counter[8] ),
    .A2(_2116_),
    .B(\soc.spi_video_ram_1.sram_sck_fall_edge ),
    .C(\soc.spi_video_ram_1.current_state[4] ),
    .ZN(_2117_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4710_ (.I0(net9),
    .I1(\soc.spi_video_ram_1.read_value[0] ),
    .S(_2117_),
    .Z(_2118_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4711_ (.I(_2118_),
    .Z(_0189_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4712_ (.A1(net10),
    .A2(_2117_),
    .ZN(_2119_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4713_ (.A1(_1349_),
    .A2(_2117_),
    .B(_2119_),
    .ZN(_0190_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4714_ (.I0(net11),
    .I1(\soc.spi_video_ram_1.read_value[2] ),
    .S(_2117_),
    .Z(_2120_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4715_ (.I(_2120_),
    .Z(_0191_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4716_ (.I0(net12),
    .I1(\soc.spi_video_ram_1.read_value[3] ),
    .S(_2117_),
    .Z(_2121_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4717_ (.I(_2121_),
    .Z(_0192_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4718_ (.I(_1670_),
    .Z(_2122_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4719_ (.I(_1482_),
    .ZN(_2123_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _4720_ (.A1(_1412_),
    .A2(_1420_),
    .A3(_1440_),
    .B(_2123_),
    .ZN(_2124_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4721_ (.I(_2124_),
    .Z(_2125_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4722_ (.A1(\soc.rom_encoder_0.output_buffer[1] ),
    .A2(_2125_),
    .ZN(_2126_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4723_ (.A1(\soc.rom_encoder_0.output_buffer[5] ),
    .A2(_1670_),
    .B1(_1672_),
    .B2(\soc.rom_encoder_0.request_address[4] ),
    .ZN(_2127_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4724_ (.A1(_2122_),
    .A2(_2126_),
    .B(_2127_),
    .ZN(_0193_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4725_ (.A1(\soc.rom_encoder_0.output_buffer[2] ),
    .A2(_2125_),
    .ZN(_2128_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4726_ (.A1(\soc.rom_encoder_0.output_buffer[6] ),
    .A2(_1670_),
    .B1(_1672_),
    .B2(\soc.rom_encoder_0.request_address[5] ),
    .ZN(_2129_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4727_ (.A1(_2122_),
    .A2(_2128_),
    .B(_2129_),
    .ZN(_0194_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4728_ (.A1(\soc.rom_encoder_0.output_buffer[3] ),
    .A2(_2125_),
    .ZN(_2130_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4729_ (.A1(\soc.rom_encoder_0.output_buffer[7] ),
    .A2(_1670_),
    .ZN(_2131_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4730_ (.A1(\soc.rom_encoder_0.request_address[6] ),
    .A2(_1672_),
    .ZN(_2132_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4731_ (.A1(_1671_),
    .A2(_2130_),
    .B(_2131_),
    .C(_2132_),
    .ZN(_0195_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4732_ (.A1(\soc.rom_encoder_0.request_data_out[0] ),
    .A2(_1481_),
    .Z(_2133_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _4733_ (.A1(\soc.rom_encoder_0.request_address[7] ),
    .A2(_1650_),
    .B1(_2125_),
    .B2(\soc.rom_encoder_0.output_buffer[4] ),
    .C(_2133_),
    .ZN(_2134_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4734_ (.A1(\soc.rom_encoder_0.output_buffer[8] ),
    .A2(_1671_),
    .ZN(_2135_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4735_ (.A1(_2122_),
    .A2(_2134_),
    .B(_2135_),
    .ZN(_0196_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4736_ (.A1(\soc.rom_encoder_0.request_data_out[1] ),
    .A2(_1481_),
    .Z(_2136_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _4737_ (.A1(\soc.rom_encoder_0.request_address[8] ),
    .A2(_1650_),
    .B1(_2125_),
    .B2(\soc.rom_encoder_0.output_buffer[5] ),
    .C(_2136_),
    .ZN(_2137_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4738_ (.I(_1670_),
    .Z(_2138_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4739_ (.A1(\soc.rom_encoder_0.output_buffer[9] ),
    .A2(_2138_),
    .ZN(_2139_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4740_ (.A1(_2122_),
    .A2(_2137_),
    .B(_2139_),
    .ZN(_0197_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4741_ (.A1(\soc.rom_encoder_0.request_data_out[2] ),
    .A2(_1481_),
    .Z(_2140_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _4742_ (.A1(\soc.rom_encoder_0.request_address[9] ),
    .A2(_1650_),
    .B1(_2125_),
    .B2(\soc.rom_encoder_0.output_buffer[6] ),
    .C(_2140_),
    .ZN(_2141_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4743_ (.A1(\soc.rom_encoder_0.output_buffer[10] ),
    .A2(_2138_),
    .ZN(_2142_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4744_ (.A1(_2122_),
    .A2(_2141_),
    .B(_2142_),
    .ZN(_0198_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4745_ (.A1(\soc.rom_encoder_0.request_data_out[3] ),
    .A2(_1481_),
    .Z(_2143_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _4746_ (.A1(\soc.rom_encoder_0.request_address[10] ),
    .A2(_1650_),
    .B1(_2125_),
    .B2(\soc.rom_encoder_0.output_buffer[7] ),
    .C(_2143_),
    .ZN(_2144_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4747_ (.A1(\soc.rom_encoder_0.output_buffer[11] ),
    .A2(_2138_),
    .ZN(_2145_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4748_ (.A1(_2122_),
    .A2(_2144_),
    .B(_2145_),
    .ZN(_0199_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4749_ (.A1(\soc.rom_encoder_0.request_data_out[4] ),
    .A2(_1481_),
    .Z(_2146_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _4750_ (.A1(\soc.rom_encoder_0.request_address[11] ),
    .A2(_1650_),
    .B1(_2125_),
    .B2(\soc.rom_encoder_0.output_buffer[8] ),
    .C(_2146_),
    .ZN(_2147_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4751_ (.A1(\soc.rom_encoder_0.output_buffer[12] ),
    .A2(_2138_),
    .ZN(_2148_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4752_ (.A1(_2122_),
    .A2(_2147_),
    .B(_2148_),
    .ZN(_0200_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4753_ (.A1(\soc.rom_encoder_0.request_data_out[5] ),
    .A2(_1481_),
    .Z(_2149_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _4754_ (.A1(\soc.rom_encoder_0.request_address[12] ),
    .A2(_1650_),
    .B1(_2125_),
    .B2(\soc.rom_encoder_0.output_buffer[9] ),
    .C(_2149_),
    .ZN(_2150_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4755_ (.A1(\soc.rom_encoder_0.output_buffer[13] ),
    .A2(_2138_),
    .ZN(_2151_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4756_ (.A1(_2122_),
    .A2(_2150_),
    .B(_2151_),
    .ZN(_0201_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4757_ (.A1(\soc.rom_encoder_0.request_data_out[6] ),
    .A2(_1481_),
    .Z(_2152_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _4758_ (.A1(\soc.rom_encoder_0.request_address[13] ),
    .A2(_1650_),
    .B1(_2125_),
    .B2(\soc.rom_encoder_0.output_buffer[10] ),
    .C(_2152_),
    .ZN(_2153_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4759_ (.A1(\soc.rom_encoder_0.output_buffer[14] ),
    .A2(_2138_),
    .ZN(_2154_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4760_ (.A1(_2122_),
    .A2(_2153_),
    .B(_2154_),
    .ZN(_0202_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4761_ (.A1(\soc.rom_encoder_0.request_data_out[7] ),
    .A2(_1481_),
    .Z(_2155_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _4762_ (.A1(\soc.rom_encoder_0.request_address[14] ),
    .A2(_1650_),
    .B1(_2124_),
    .B2(\soc.rom_encoder_0.output_buffer[11] ),
    .C(_2155_),
    .ZN(_2156_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4763_ (.A1(\soc.rom_encoder_0.output_buffer[15] ),
    .A2(_2138_),
    .ZN(_2157_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4764_ (.A1(_2122_),
    .A2(_2156_),
    .B(_2157_),
    .ZN(_0203_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4765_ (.A1(_1437_),
    .A2(_1482_),
    .B(\soc.rom_encoder_0.output_buffer[12] ),
    .ZN(_2158_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4766_ (.A1(\soc.rom_encoder_0.request_data_out[8] ),
    .A2(_1481_),
    .ZN(_2159_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4767_ (.A1(\soc.rom_encoder_0.request_write ),
    .A2(_1656_),
    .B(_2158_),
    .C(_2159_),
    .ZN(_2160_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4768_ (.A1(_1441_),
    .A2(_2160_),
    .ZN(_2161_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4769_ (.A1(\soc.rom_encoder_0.output_buffer[16] ),
    .A2(_2138_),
    .ZN(_2162_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4770_ (.A1(_1671_),
    .A2(_2161_),
    .B(_2162_),
    .ZN(_0204_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4771_ (.A1(_1421_),
    .A2(_1442_),
    .ZN(_2163_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4772_ (.A1(\soc.rom_encoder_0.request_data_out[9] ),
    .A2(_1434_),
    .ZN(_2164_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4773_ (.A1(\soc.rom_encoder_0.current_state[1] ),
    .A2(_2164_),
    .ZN(_2165_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _4774_ (.A1(\soc.rom_encoder_0.output_buffer[13] ),
    .A2(_2163_),
    .B1(_2165_),
    .B2(_1435_),
    .C(_1441_),
    .ZN(_2166_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4775_ (.A1(\soc.rom_encoder_0.output_buffer[17] ),
    .A2(_2138_),
    .ZN(_2167_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4776_ (.A1(_1671_),
    .A2(_2166_),
    .B(_2167_),
    .ZN(_0205_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4777_ (.A1(\soc.rom_encoder_0.output_buffer[14] ),
    .A2(_1417_),
    .B1(_1442_),
    .B2(\soc.rom_encoder_0.request_data_out[10] ),
    .ZN(_2168_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4778_ (.A1(_1413_),
    .A2(_2168_),
    .ZN(_2169_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _4779_ (.A1(\soc.rom_encoder_0.output_buffer[14] ),
    .A2(_1436_),
    .B(_2169_),
    .C(_1441_),
    .ZN(_2170_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4780_ (.A1(\soc.rom_encoder_0.output_buffer[18] ),
    .A2(_2138_),
    .ZN(_2171_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4781_ (.A1(_1671_),
    .A2(_2170_),
    .B(_2171_),
    .ZN(_0206_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4782_ (.A1(\soc.rom_encoder_0.output_buffer[15] ),
    .A2(_1417_),
    .B1(_1442_),
    .B2(\soc.rom_encoder_0.request_data_out[11] ),
    .ZN(_2172_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4783_ (.A1(_1413_),
    .A2(_2172_),
    .ZN(_2173_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _4784_ (.A1(\soc.rom_encoder_0.output_buffer[15] ),
    .A2(_1436_),
    .B(_2173_),
    .C(_1441_),
    .ZN(_2174_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4785_ (.A1(\soc.rom_encoder_0.output_buffer[19] ),
    .A2(_1670_),
    .ZN(_2175_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4786_ (.A1(_1671_),
    .A2(_2174_),
    .B(_2175_),
    .ZN(_0207_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4787_ (.A1(_0674_),
    .A2(\soc.spi_video_ram_1.sram_sck_rise_edge ),
    .Z(_2176_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4788_ (.A1(_0720_),
    .A2(_2176_),
    .ZN(_2177_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4789_ (.A1(_0776_),
    .A2(_2177_),
    .Z(_2178_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4790_ (.A1(_0776_),
    .A2(_2177_),
    .ZN(_2179_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _4791_ (.A1(\soc.spi_video_ram_1.state_sram_clk_counter[0] ),
    .A2(_0684_),
    .A3(_0715_),
    .ZN(_2180_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _4792_ (.A1(_2180_),
    .A2(_0704_),
    .B1(_0721_),
    .B2(_0703_),
    .C(_1575_),
    .ZN(_2181_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _4793_ (.A1(_0689_),
    .A2(_0705_),
    .A3(_2181_),
    .Z(_2182_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4794_ (.A1(_2178_),
    .A2(_2179_),
    .A3(_2182_),
    .ZN(_0208_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4795_ (.A1(_0758_),
    .A2(_2178_),
    .ZN(_2183_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4796_ (.A1(_0764_),
    .A2(_2177_),
    .B(_2182_),
    .C(_2183_),
    .ZN(_0209_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4797_ (.A1(\soc.spi_video_ram_1.current_state[3] ),
    .A2(_0764_),
    .ZN(_2184_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4798_ (.A1(_0810_),
    .A2(_2176_),
    .A3(_2184_),
    .ZN(_2185_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4799_ (.A1(_2176_),
    .A2(_2184_),
    .ZN(_2186_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4800_ (.A1(_0759_),
    .A2(_2186_),
    .ZN(_2187_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4801_ (.A1(_2182_),
    .A2(_2185_),
    .A3(_2187_),
    .ZN(_0210_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4802_ (.A1(_0752_),
    .A2(_2185_),
    .Z(_2188_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4803_ (.A1(_1796_),
    .A2(_2188_),
    .ZN(_0211_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4804_ (.A1(_0720_),
    .A2(_1383_),
    .ZN(_2189_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4805_ (.A1(_0720_),
    .A2(_0754_),
    .B(_2176_),
    .C(_2189_),
    .ZN(_2190_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4806_ (.A1(_0749_),
    .A2(_2176_),
    .B(_2182_),
    .C(_2190_),
    .ZN(_0212_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _4807_ (.A1(_0749_),
    .A2(_0753_),
    .A3(_2176_),
    .A4(_2184_),
    .ZN(_2191_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4808_ (.A1(\soc.spi_video_ram_1.buffer_index[5] ),
    .A2(_2191_),
    .Z(_2192_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4809_ (.A1(_1796_),
    .A2(_2192_),
    .ZN(_0213_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4810_ (.A1(\soc.spi_video_ram_1.state_sram_clk_counter[8] ),
    .A2(_2116_),
    .B(_0729_),
    .ZN(_0214_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4811_ (.I0(\soc.spi_video_ram_1.fifo_in_address[0] ),
    .I1(\soc.cpu.AReg.data[0] ),
    .S(_2018_),
    .Z(_2193_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4812_ (.I(_2193_),
    .Z(_0215_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4813_ (.I0(\soc.spi_video_ram_1.fifo_in_address[1] ),
    .I1(\soc.cpu.AReg.data[1] ),
    .S(_2018_),
    .Z(_2194_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4814_ (.I(_2194_),
    .Z(_0216_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4815_ (.I0(\soc.spi_video_ram_1.fifo_in_address[2] ),
    .I1(\soc.cpu.AReg.data[2] ),
    .S(_2018_),
    .Z(_2195_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4816_ (.I(_2195_),
    .Z(_0217_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4817_ (.I0(\soc.spi_video_ram_1.fifo_in_address[3] ),
    .I1(\soc.cpu.AReg.data[3] ),
    .S(_2018_),
    .Z(_2196_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4818_ (.I(_2196_),
    .Z(_0218_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4819_ (.I0(\soc.spi_video_ram_1.fifo_in_address[4] ),
    .I1(\soc.cpu.AReg.data[4] ),
    .S(_2018_),
    .Z(_2197_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4820_ (.I(_2197_),
    .Z(_0219_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4821_ (.I0(\soc.spi_video_ram_1.fifo_in_address[5] ),
    .I1(\soc.cpu.AReg.data[5] ),
    .S(_2018_),
    .Z(_2198_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4822_ (.I(_2198_),
    .Z(_0220_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4823_ (.I0(\soc.spi_video_ram_1.fifo_in_address[6] ),
    .I1(\soc.cpu.AReg.data[6] ),
    .S(_2018_),
    .Z(_2199_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4824_ (.I(_2199_),
    .Z(_0221_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4825_ (.I0(\soc.spi_video_ram_1.fifo_in_address[7] ),
    .I1(\soc.cpu.AReg.data[7] ),
    .S(_0748_),
    .Z(_2200_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4826_ (.I(_2200_),
    .Z(_0222_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4827_ (.I0(\soc.spi_video_ram_1.fifo_in_address[8] ),
    .I1(\soc.cpu.AReg.data[8] ),
    .S(_0748_),
    .Z(_2201_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4828_ (.I(_2201_),
    .Z(_0223_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4829_ (.I0(\soc.spi_video_ram_1.fifo_in_address[9] ),
    .I1(\soc.cpu.AReg.data[9] ),
    .S(_0748_),
    .Z(_2202_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4830_ (.I(_2202_),
    .Z(_0224_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4831_ (.I0(\soc.spi_video_ram_1.fifo_in_address[10] ),
    .I1(\soc.cpu.AReg.data[10] ),
    .S(_0748_),
    .Z(_2203_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4832_ (.I(_2203_),
    .Z(_0225_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4833_ (.I0(\soc.spi_video_ram_1.fifo_in_address[11] ),
    .I1(\soc.cpu.AReg.data[11] ),
    .S(_0748_),
    .Z(_2204_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4834_ (.I(_2204_),
    .Z(_0226_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4835_ (.I0(\soc.spi_video_ram_1.fifo_in_address[12] ),
    .I1(\soc.cpu.AReg.data[12] ),
    .S(_0748_),
    .Z(_2205_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4836_ (.I(_2205_),
    .Z(_0227_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4837_ (.A1(\soc.video_generator_1.h_count[4] ),
    .A2(_1132_),
    .ZN(_2206_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _4838_ (.A1(_1216_),
    .A2(_1131_),
    .A3(_2206_),
    .ZN(_2207_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _4839_ (.A1(\soc.spi_video_ram_1.initialized ),
    .A2(\soc.video_generator_1.h_count[1] ),
    .A3(_1189_),
    .A4(_2207_),
    .ZN(_2208_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _4840_ (.A1(_1356_),
    .A2(_1455_),
    .A3(_2208_),
    .B(_0705_),
    .ZN(_2209_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4841_ (.A1(\soc.spi_video_ram_1.start_read ),
    .A2(_0705_),
    .B(_2209_),
    .ZN(_2210_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4842_ (.A1(_0691_),
    .A2(_2210_),
    .ZN(_0228_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4843_ (.A1(_0727_),
    .A2(_0722_),
    .B(_0691_),
    .ZN(_0229_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4844_ (.I(\soc.spi_video_ram_1.fifo_write_request ),
    .ZN(_2211_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4845_ (.A1(_1949_),
    .A2(_0740_),
    .B(_2211_),
    .ZN(_2212_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4846_ (.A1(_0698_),
    .A2(_2212_),
    .Z(_2213_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4847_ (.A1(_0698_),
    .A2(_2212_),
    .B(_1955_),
    .ZN(_2214_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4848_ (.A1(_2213_),
    .A2(_2214_),
    .ZN(_0230_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4849_ (.A1(_0694_),
    .A2(_2213_),
    .B(_1955_),
    .ZN(_2215_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4850_ (.A1(_0694_),
    .A2(_2213_),
    .B(_2215_),
    .ZN(_0231_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _4851_ (.A1(\soc.spi_video_ram_1.write_fifo.write_pointer[2] ),
    .A2(_0738_),
    .ZN(_2216_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _4852_ (.I(_2216_),
    .Z(_2217_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4853_ (.A1(_0694_),
    .A2(_2213_),
    .B(_0700_),
    .ZN(_2218_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4854_ (.A1(_2212_),
    .A2(_2217_),
    .B(_2218_),
    .ZN(_2219_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4855_ (.A1(_0691_),
    .A2(_2219_),
    .ZN(_0232_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _4856_ (.A1(_1461_),
    .A2(_1951_),
    .A3(_1952_),
    .ZN(_0233_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _4857_ (.A1(_1461_),
    .A2(_1953_),
    .A3(_1954_),
    .ZN(_0234_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4858_ (.A1(_1955_),
    .A2(_1956_),
    .Z(_2220_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4859_ (.I(_2220_),
    .Z(_0235_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4860_ (.A1(\soc.rom_encoder_0.current_state[1] ),
    .A2(_1406_),
    .ZN(_2221_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4861_ (.A1(_1426_),
    .A2(_2221_),
    .ZN(_2222_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _4862_ (.A1(_1407_),
    .A2(_1422_),
    .ZN(_2223_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4863_ (.A1(\soc.rom_encoder_0.current_state[1] ),
    .A2(_1406_),
    .ZN(_2224_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4864_ (.A1(_1426_),
    .A2(_2224_),
    .ZN(_2225_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4865_ (.I(\soc.rom_encoder_0.input_bits_left[3] ),
    .ZN(_2226_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4866_ (.I(\soc.rom_encoder_0.input_bits_left[4] ),
    .ZN(_2227_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4867_ (.A1(\soc.rom_encoder_0.input_bits_left[2] ),
    .A2(_2226_),
    .A3(_2227_),
    .ZN(_2228_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4868_ (.A1(\soc.rom_encoder_0.request_write ),
    .A2(_1417_),
    .B(_2222_),
    .ZN(_2229_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4869_ (.A1(_2225_),
    .A2(_2228_),
    .B(_1403_),
    .C(_2229_),
    .ZN(_2230_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4870_ (.A1(net18),
    .A2(_2230_),
    .ZN(_2231_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4871_ (.A1(_2222_),
    .A2(_2223_),
    .B(_2231_),
    .ZN(_2232_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4872_ (.A1(\soc.rom_encoder_0.input_bits_left[2] ),
    .A2(_2232_),
    .ZN(_2233_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4873_ (.A1(\soc.rom_encoder_0.input_bits_left[2] ),
    .A2(_2232_),
    .ZN(_2234_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4874_ (.A1(_1426_),
    .A2(_2234_),
    .ZN(_2235_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4875_ (.A1(_2233_),
    .A2(_2235_),
    .ZN(_0236_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4876_ (.A1(_2222_),
    .A2(_2231_),
    .ZN(_2236_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4877_ (.A1(_2226_),
    .A2(_2234_),
    .ZN(_2237_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4878_ (.A1(\soc.rom_encoder_0.input_bits_left[2] ),
    .A2(_2232_),
    .B(\soc.rom_encoder_0.input_bits_left[3] ),
    .ZN(_2238_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4879_ (.A1(_2236_),
    .A2(_2237_),
    .A3(_2238_),
    .ZN(_0237_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4880_ (.A1(\soc.rom_encoder_0.input_bits_left[4] ),
    .A2(_2237_),
    .Z(_2239_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4881_ (.A1(_2236_),
    .A2(_2239_),
    .ZN(_0238_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4882_ (.I(\soc.rom_encoder_0.input_buffer[0] ),
    .ZN(_2240_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4883_ (.A1(_1403_),
    .A2(_2223_),
    .ZN(_2241_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4884_ (.I(_2241_),
    .Z(_2242_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4885_ (.I(_2241_),
    .Z(_2243_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4886_ (.A1(net5),
    .A2(_2243_),
    .B(_1955_),
    .ZN(_2244_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4887_ (.A1(_2240_),
    .A2(_2242_),
    .B(_2244_),
    .ZN(_0239_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4888_ (.I(\soc.rom_encoder_0.input_buffer[1] ),
    .ZN(_2245_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4889_ (.A1(net6),
    .A2(_2243_),
    .B(_1955_),
    .ZN(_2246_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4890_ (.A1(_2245_),
    .A2(_2242_),
    .B(_2246_),
    .ZN(_0240_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4891_ (.I(\soc.rom_encoder_0.input_buffer[2] ),
    .ZN(_2247_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4892_ (.A1(net7),
    .A2(_2243_),
    .B(_1955_),
    .ZN(_2248_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4893_ (.A1(_2247_),
    .A2(_2242_),
    .B(_2248_),
    .ZN(_0241_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4894_ (.I(\soc.rom_encoder_0.input_buffer[3] ),
    .ZN(_2249_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4895_ (.I(_0675_),
    .Z(_2250_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4896_ (.A1(net8),
    .A2(_2243_),
    .B(_2250_),
    .ZN(_2251_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4897_ (.A1(_2249_),
    .A2(_2242_),
    .B(_2251_),
    .ZN(_0242_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4898_ (.I(\soc.rom_encoder_0.input_buffer[4] ),
    .ZN(_2252_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4899_ (.A1(\soc.rom_encoder_0.input_buffer[0] ),
    .A2(_2243_),
    .B(_2250_),
    .ZN(_2253_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4900_ (.A1(_2252_),
    .A2(_2242_),
    .B(_2253_),
    .ZN(_0243_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4901_ (.I(\soc.rom_encoder_0.input_buffer[5] ),
    .ZN(_2254_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4902_ (.A1(\soc.rom_encoder_0.input_buffer[1] ),
    .A2(_2243_),
    .B(_2250_),
    .ZN(_2255_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4903_ (.A1(_2254_),
    .A2(_2242_),
    .B(_2255_),
    .ZN(_0244_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4904_ (.I(\soc.rom_encoder_0.input_buffer[6] ),
    .ZN(_2256_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4905_ (.A1(\soc.rom_encoder_0.input_buffer[2] ),
    .A2(_2243_),
    .B(_2250_),
    .ZN(_2257_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4906_ (.A1(_2256_),
    .A2(_2242_),
    .B(_2257_),
    .ZN(_0245_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4907_ (.I(\soc.rom_encoder_0.input_buffer[7] ),
    .ZN(_2258_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4908_ (.A1(\soc.rom_encoder_0.input_buffer[3] ),
    .A2(_2243_),
    .B(_2250_),
    .ZN(_2259_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4909_ (.A1(_2258_),
    .A2(_2242_),
    .B(_2259_),
    .ZN(_0246_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4910_ (.I(\soc.rom_encoder_0.input_buffer[8] ),
    .ZN(_2260_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4911_ (.A1(\soc.rom_encoder_0.input_buffer[4] ),
    .A2(_2241_),
    .B(_2250_),
    .ZN(_2261_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4912_ (.A1(_2260_),
    .A2(_2242_),
    .B(_2261_),
    .ZN(_0247_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4913_ (.I(\soc.rom_encoder_0.input_buffer[9] ),
    .ZN(_2262_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4914_ (.A1(\soc.rom_encoder_0.input_buffer[5] ),
    .A2(_2241_),
    .B(_2250_),
    .ZN(_2263_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4915_ (.A1(_2262_),
    .A2(_2242_),
    .B(_2263_),
    .ZN(_0248_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4916_ (.I(\soc.rom_encoder_0.input_buffer[10] ),
    .ZN(_2264_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4917_ (.A1(\soc.rom_encoder_0.input_buffer[6] ),
    .A2(_2241_),
    .B(_2250_),
    .ZN(_2265_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4918_ (.A1(_2264_),
    .A2(_2243_),
    .B(_2265_),
    .ZN(_0249_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4919_ (.I(\soc.rom_encoder_0.input_buffer[11] ),
    .ZN(_2266_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4920_ (.A1(\soc.rom_encoder_0.input_buffer[7] ),
    .A2(_2241_),
    .B(_2250_),
    .ZN(_2267_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4921_ (.A1(_2266_),
    .A2(_2243_),
    .B(_2267_),
    .ZN(_0250_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4922_ (.A1(\soc.rom_encoder_0.current_state[2] ),
    .A2(_1422_),
    .ZN(_2268_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4923_ (.I0(\soc.hack_rom_request ),
    .I1(\soc.rom_loader.rom_request ),
    .S(\soc.rom_encoder_0.write_enable ),
    .Z(_2269_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _4924_ (.A1(_1403_),
    .A2(_0674_),
    .A3(_2268_),
    .A4(_2269_),
    .ZN(_2270_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 _4925_ (.I(_2270_),
    .Z(_2271_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _4926_ (.I(_2271_),
    .Z(_2272_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4927_ (.A1(\soc.rom_encoder_0.request_write ),
    .A2(_2272_),
    .ZN(_2273_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4928_ (.A1(_2089_),
    .A2(_2272_),
    .B(_2273_),
    .ZN(_0251_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4929_ (.I0(\soc.rom_encoder_0.data_out[0] ),
    .I1(\soc.rom_encoder_0.request_data_out[0] ),
    .S(_2272_),
    .Z(_2274_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4930_ (.I(_2274_),
    .Z(_0252_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4931_ (.I0(\soc.rom_encoder_0.data_out[1] ),
    .I1(\soc.rom_encoder_0.request_data_out[1] ),
    .S(_2272_),
    .Z(_2275_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4932_ (.I(_2275_),
    .Z(_0253_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _4933_ (.I(_2271_),
    .Z(_2276_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4934_ (.I0(\soc.rom_encoder_0.data_out[2] ),
    .I1(\soc.rom_encoder_0.request_data_out[2] ),
    .S(_2276_),
    .Z(_2277_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4935_ (.I(_2277_),
    .Z(_0254_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4936_ (.I0(\soc.rom_encoder_0.data_out[3] ),
    .I1(\soc.rom_encoder_0.request_data_out[3] ),
    .S(_2276_),
    .Z(_2278_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4937_ (.I(_2278_),
    .Z(_0255_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4938_ (.I0(\soc.rom_encoder_0.data_out[4] ),
    .I1(\soc.rom_encoder_0.request_data_out[4] ),
    .S(_2276_),
    .Z(_2279_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4939_ (.I(_2279_),
    .Z(_0256_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4940_ (.I0(\soc.rom_encoder_0.data_out[5] ),
    .I1(\soc.rom_encoder_0.request_data_out[5] ),
    .S(_2276_),
    .Z(_2280_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4941_ (.I(_2280_),
    .Z(_0257_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4942_ (.I0(\soc.rom_encoder_0.data_out[6] ),
    .I1(\soc.rom_encoder_0.request_data_out[6] ),
    .S(_2276_),
    .Z(_2281_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4943_ (.I(_2281_),
    .Z(_0258_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4944_ (.I0(\soc.rom_encoder_0.data_out[7] ),
    .I1(\soc.rom_encoder_0.request_data_out[7] ),
    .S(_2276_),
    .Z(_2282_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4945_ (.I(_2282_),
    .Z(_0259_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4946_ (.I0(\soc.rom_encoder_0.data_out[8] ),
    .I1(\soc.rom_encoder_0.request_data_out[8] ),
    .S(_2276_),
    .Z(_2283_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4947_ (.I(_2283_),
    .Z(_0260_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4948_ (.I0(\soc.rom_encoder_0.data_out[9] ),
    .I1(\soc.rom_encoder_0.request_data_out[9] ),
    .S(_2276_),
    .Z(_2284_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4949_ (.I(_2284_),
    .Z(_0261_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4950_ (.I0(\soc.rom_encoder_0.data_out[10] ),
    .I1(\soc.rom_encoder_0.request_data_out[10] ),
    .S(_2276_),
    .Z(_2285_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4951_ (.I(_2285_),
    .Z(_0262_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4952_ (.I0(\soc.rom_encoder_0.data_out[11] ),
    .I1(\soc.rom_encoder_0.request_data_out[11] ),
    .S(_2276_),
    .Z(_2286_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4953_ (.I(_2286_),
    .Z(_0263_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _4954_ (.I(_2271_),
    .Z(_2287_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4955_ (.I0(\soc.rom_encoder_0.data_out[12] ),
    .I1(\soc.rom_encoder_0.request_data_out[12] ),
    .S(_2287_),
    .Z(_2288_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4956_ (.I(_2288_),
    .Z(_0264_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4957_ (.I0(\soc.rom_encoder_0.data_out[13] ),
    .I1(\soc.rom_encoder_0.request_data_out[13] ),
    .S(_2287_),
    .Z(_2289_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4958_ (.I(_2289_),
    .Z(_0265_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4959_ (.I0(\soc.rom_encoder_0.data_out[14] ),
    .I1(\soc.rom_encoder_0.request_data_out[14] ),
    .S(_2287_),
    .Z(_2290_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4960_ (.I(_2290_),
    .Z(_0266_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4961_ (.I0(\soc.rom_encoder_0.data_out[15] ),
    .I1(\soc.rom_encoder_0.request_data_out[15] ),
    .S(_2287_),
    .Z(_2291_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4962_ (.I(_2291_),
    .Z(_0267_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _4963_ (.I(\soc.rom_encoder_0.write_enable ),
    .Z(_2292_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _4964_ (.I(_2292_),
    .Z(_2293_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4965_ (.I0(\soc.cpu.PC.REG.data[0] ),
    .I1(\soc.rom_loader.current_address[0] ),
    .S(_2293_),
    .Z(_2294_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4966_ (.I0(_2294_),
    .I1(\soc.rom_encoder_0.request_address[0] ),
    .S(_2287_),
    .Z(_2295_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4967_ (.I(_2295_),
    .Z(_0268_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4968_ (.I0(\soc.cpu.PC.REG.data[1] ),
    .I1(\soc.rom_loader.current_address[1] ),
    .S(_2293_),
    .Z(_2296_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4969_ (.I0(_2296_),
    .I1(\soc.rom_encoder_0.request_address[1] ),
    .S(_2287_),
    .Z(_2297_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4970_ (.I(_2297_),
    .Z(_0269_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4971_ (.I0(\soc.cpu.PC.REG.data[2] ),
    .I1(\soc.rom_loader.current_address[2] ),
    .S(_2293_),
    .Z(_2298_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4972_ (.I0(_2298_),
    .I1(\soc.rom_encoder_0.request_address[2] ),
    .S(_2287_),
    .Z(_2299_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4973_ (.I(_2299_),
    .Z(_0270_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4974_ (.I(\soc.cpu.PC.REG.data[3] ),
    .ZN(_2300_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4975_ (.A1(_2293_),
    .A2(_2300_),
    .ZN(_2301_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4976_ (.A1(_2293_),
    .A2(\soc.rom_loader.current_address[3] ),
    .B(_2301_),
    .ZN(_2302_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4977_ (.A1(\soc.rom_encoder_0.request_address[3] ),
    .A2(_2272_),
    .ZN(_2303_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4978_ (.A1(_2272_),
    .A2(_2302_),
    .B(_2303_),
    .ZN(_0271_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4979_ (.I0(\soc.cpu.PC.REG.data[4] ),
    .I1(\soc.rom_loader.current_address[4] ),
    .S(_2292_),
    .Z(_2304_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4980_ (.I0(_2304_),
    .I1(\soc.rom_encoder_0.request_address[4] ),
    .S(_2287_),
    .Z(_2305_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4981_ (.I(_2305_),
    .Z(_0272_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4982_ (.I0(\soc.cpu.PC.REG.data[5] ),
    .I1(\soc.rom_loader.current_address[5] ),
    .S(_2292_),
    .Z(_2306_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4983_ (.I0(_2306_),
    .I1(\soc.rom_encoder_0.request_address[5] ),
    .S(_2287_),
    .Z(_2307_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4984_ (.I(_2307_),
    .Z(_0273_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4985_ (.I0(\soc.cpu.PC.REG.data[6] ),
    .I1(\soc.rom_loader.current_address[6] ),
    .S(_2292_),
    .Z(_2308_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4986_ (.I0(_2308_),
    .I1(\soc.rom_encoder_0.request_address[6] ),
    .S(_2287_),
    .Z(_2309_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4987_ (.I(_2309_),
    .Z(_0274_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4988_ (.I(\soc.cpu.PC.REG.data[7] ),
    .ZN(_2310_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4989_ (.A1(_2293_),
    .A2(_2310_),
    .ZN(_2311_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4990_ (.A1(_2293_),
    .A2(\soc.rom_loader.current_address[7] ),
    .B(_2311_),
    .ZN(_2312_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4991_ (.A1(\soc.rom_encoder_0.request_address[7] ),
    .A2(_2272_),
    .ZN(_2313_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4992_ (.A1(_2272_),
    .A2(_2312_),
    .B(_2313_),
    .ZN(_0275_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4993_ (.I0(\soc.cpu.PC.REG.data[8] ),
    .I1(\soc.rom_loader.current_address[8] ),
    .S(_2292_),
    .Z(_2314_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4994_ (.I0(_2314_),
    .I1(\soc.rom_encoder_0.request_address[8] ),
    .S(_2271_),
    .Z(_2315_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4995_ (.I(_2315_),
    .Z(_0276_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4996_ (.I0(\soc.cpu.PC.REG.data[9] ),
    .I1(\soc.rom_loader.current_address[9] ),
    .S(_2292_),
    .Z(_2316_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4997_ (.I0(_2316_),
    .I1(\soc.rom_encoder_0.request_address[9] ),
    .S(_2271_),
    .Z(_2317_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4998_ (.I(_2317_),
    .Z(_0277_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4999_ (.I(\soc.cpu.PC.REG.data[10] ),
    .ZN(_2318_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5000_ (.A1(_2293_),
    .A2(_2318_),
    .ZN(_2319_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5001_ (.A1(_2293_),
    .A2(\soc.rom_loader.current_address[10] ),
    .B(_2319_),
    .ZN(_2320_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5002_ (.A1(\soc.rom_encoder_0.request_address[10] ),
    .A2(_2272_),
    .ZN(_2321_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5003_ (.A1(_2272_),
    .A2(_2320_),
    .B(_2321_),
    .ZN(_0278_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5004_ (.I0(\soc.cpu.PC.REG.data[11] ),
    .I1(\soc.rom_loader.current_address[11] ),
    .S(_2292_),
    .Z(_2322_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5005_ (.I0(_2322_),
    .I1(\soc.rom_encoder_0.request_address[11] ),
    .S(_2271_),
    .Z(_2323_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5006_ (.I(_2323_),
    .Z(_0279_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5007_ (.I0(\soc.cpu.PC.REG.data[12] ),
    .I1(\soc.rom_loader.current_address[12] ),
    .S(_2292_),
    .Z(_2324_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5008_ (.I0(_2324_),
    .I1(\soc.rom_encoder_0.request_address[12] ),
    .S(_2271_),
    .Z(_2325_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5009_ (.I(_2325_),
    .Z(_0280_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5010_ (.I0(\soc.cpu.PC.REG.data[13] ),
    .I1(\soc.rom_loader.current_address[13] ),
    .S(_2292_),
    .Z(_2326_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5011_ (.I0(_2326_),
    .I1(\soc.rom_encoder_0.request_address[13] ),
    .S(_2271_),
    .Z(_2327_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5012_ (.I(_2327_),
    .Z(_0281_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5013_ (.I0(\soc.cpu.PC.REG.data[14] ),
    .I1(\soc.rom_loader.current_address[14] ),
    .S(_2292_),
    .Z(_2328_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5014_ (.I0(_2328_),
    .I1(\soc.rom_encoder_0.request_address[14] ),
    .S(_2271_),
    .Z(_2329_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5015_ (.I(_2329_),
    .Z(_0282_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5016_ (.A1(_1492_),
    .A2(_1508_),
    .ZN(_2330_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5017_ (.A1(\soc.ram_encoder_0.initializing_step[4] ),
    .A2(\soc.ram_encoder_0.initializing_step[3] ),
    .ZN(_2331_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5018_ (.A1(_2331_),
    .A2(_1508_),
    .ZN(_2332_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5019_ (.A1(net58),
    .A2(_2330_),
    .A3(_2332_),
    .ZN(_2333_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5020_ (.A1(_1493_),
    .A2(\soc.ram_encoder_0.current_state[1] ),
    .ZN(_2334_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5021_ (.A1(_1488_),
    .A2(_2334_),
    .ZN(_2335_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5022_ (.A1(_2335_),
    .A2(_1516_),
    .B1(_1529_),
    .B2(\soc.ram_encoder_0.request_data_out[12] ),
    .ZN(_2336_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5023_ (.A1(_1489_),
    .A2(_1512_),
    .B(_1518_),
    .ZN(_2337_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5024_ (.A1(\soc.ram_encoder_0.initializing_step[1] ),
    .A2(\soc.ram_encoder_0.initializing_step[0] ),
    .B(_2331_),
    .C(\soc.ram_encoder_0.initializing_step[2] ),
    .ZN(_2338_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5025_ (.A1(_1492_),
    .A2(_1494_),
    .ZN(_2339_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5026_ (.A1(\soc.ram_encoder_0.output_buffer[16] ),
    .A2(_2337_),
    .B1(_2338_),
    .B2(_2339_),
    .ZN(_2340_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5027_ (.A1(_2330_),
    .A2(_2332_),
    .B1(_2336_),
    .B2(_2340_),
    .ZN(_2341_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5028_ (.A1(_0690_),
    .A2(_2341_),
    .ZN(_2342_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5029_ (.A1(_2333_),
    .A2(_2342_),
    .ZN(_0283_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _5030_ (.A1(\soc.ram_encoder_0.output_buffer[17] ),
    .A2(_1555_),
    .B1(_1529_),
    .B2(\soc.ram_encoder_0.request_data_out[13] ),
    .C(_1559_),
    .ZN(_2343_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5031_ (.A1(net59),
    .A2(_2330_),
    .ZN(_2344_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5032_ (.A1(_2330_),
    .A2(_2343_),
    .B(_2344_),
    .C(_0676_),
    .ZN(_0284_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _5033_ (.A1(\soc.ram_encoder_0.output_buffer[18] ),
    .A2(_1555_),
    .B1(_1529_),
    .B2(\soc.ram_encoder_0.request_data_out[14] ),
    .C(_1559_),
    .ZN(_2345_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5034_ (.A1(net60),
    .A2(_2330_),
    .ZN(_2346_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5035_ (.A1(_2330_),
    .A2(_2345_),
    .B(_2346_),
    .C(_0676_),
    .ZN(_0285_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _5036_ (.A1(\soc.ram_encoder_0.output_buffer[19] ),
    .A2(_1555_),
    .B1(_1529_),
    .B2(\soc.ram_encoder_0.request_data_out[15] ),
    .C(_1559_),
    .ZN(_2347_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5037_ (.A1(net61),
    .A2(_2330_),
    .ZN(_2348_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5038_ (.A1(_2330_),
    .A2(_2347_),
    .B(_2348_),
    .C(_0676_),
    .ZN(_0286_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5039_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[3][0] ),
    .I1(\soc.spi_video_ram_1.fifo_in_data[0] ),
    .S(_2217_),
    .Z(_2349_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5040_ (.I(_2349_),
    .Z(_0287_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5041_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[3][1] ),
    .I1(\soc.spi_video_ram_1.fifo_in_data[1] ),
    .S(_2217_),
    .Z(_2350_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5042_ (.I(_2350_),
    .Z(_0288_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5043_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[3][2] ),
    .I1(\soc.spi_video_ram_1.fifo_in_data[2] ),
    .S(_2217_),
    .Z(_2351_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5044_ (.I(_2351_),
    .Z(_0289_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5045_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[3][3] ),
    .I1(\soc.spi_video_ram_1.fifo_in_data[3] ),
    .S(_2217_),
    .Z(_2352_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5046_ (.I(_2352_),
    .Z(_0290_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5047_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[3][4] ),
    .I1(\soc.spi_video_ram_1.fifo_in_data[4] ),
    .S(_2217_),
    .Z(_2353_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5048_ (.I(_2353_),
    .Z(_0291_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5049_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[3][5] ),
    .I1(\soc.spi_video_ram_1.fifo_in_data[5] ),
    .S(_2217_),
    .Z(_2354_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5050_ (.I(_2354_),
    .Z(_0292_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5051_ (.A1(\soc.spi_video_ram_1.fifo_in_data[6] ),
    .A2(_2217_),
    .ZN(_2355_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5052_ (.A1(_1748_),
    .A2(_2217_),
    .B(_2355_),
    .ZN(_0293_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5053_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[3][7] ),
    .I1(\soc.spi_video_ram_1.fifo_in_data[7] ),
    .S(_2217_),
    .Z(_2356_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5054_ (.I(_2356_),
    .Z(_0294_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _5055_ (.I(_2216_),
    .Z(_2357_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5056_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[3][8] ),
    .I1(\soc.spi_video_ram_1.fifo_in_data[8] ),
    .S(_2357_),
    .Z(_2358_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5057_ (.I(_2358_),
    .Z(_0295_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5058_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[3][9] ),
    .I1(\soc.spi_video_ram_1.fifo_in_data[9] ),
    .S(_2357_),
    .Z(_2359_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5059_ (.I(_2359_),
    .Z(_0296_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5060_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[3][10] ),
    .I1(\soc.spi_video_ram_1.fifo_in_data[10] ),
    .S(_2357_),
    .Z(_2360_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5061_ (.I(_2360_),
    .Z(_0297_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5062_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[3][11] ),
    .I1(\soc.spi_video_ram_1.fifo_in_data[11] ),
    .S(_2357_),
    .Z(_2361_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5063_ (.I(_2361_),
    .Z(_0298_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5064_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[3][12] ),
    .I1(\soc.spi_video_ram_1.fifo_in_data[12] ),
    .S(_2357_),
    .Z(_2362_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5065_ (.I(_2362_),
    .Z(_0299_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5066_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[3][13] ),
    .I1(\soc.spi_video_ram_1.fifo_in_data[13] ),
    .S(_2357_),
    .Z(_2363_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5067_ (.I(_2363_),
    .Z(_0300_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5068_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[3][14] ),
    .I1(\soc.spi_video_ram_1.fifo_in_data[14] ),
    .S(_2357_),
    .Z(_2364_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5069_ (.I(_2364_),
    .Z(_0301_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5070_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[3][15] ),
    .I1(\soc.spi_video_ram_1.fifo_in_data[15] ),
    .S(_2357_),
    .Z(_2365_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5071_ (.I(_2365_),
    .Z(_0302_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5072_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[3][16] ),
    .I1(\soc.spi_video_ram_1.fifo_in_address[0] ),
    .S(_2357_),
    .Z(_2366_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5073_ (.I(_2366_),
    .Z(_0303_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5074_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[3][17] ),
    .I1(\soc.spi_video_ram_1.fifo_in_address[1] ),
    .S(_2357_),
    .Z(_2367_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5075_ (.I(_2367_),
    .Z(_0304_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _5076_ (.I(_2216_),
    .Z(_2368_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5077_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[3][18] ),
    .I1(\soc.spi_video_ram_1.fifo_in_address[2] ),
    .S(_2368_),
    .Z(_2369_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5078_ (.I(_2369_),
    .Z(_0305_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5079_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[3][19] ),
    .I1(\soc.spi_video_ram_1.fifo_in_address[3] ),
    .S(_2368_),
    .Z(_2370_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5080_ (.I(_2370_),
    .Z(_0306_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5081_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[3][20] ),
    .I1(\soc.spi_video_ram_1.fifo_in_address[4] ),
    .S(_2368_),
    .Z(_2371_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5082_ (.I(_2371_),
    .Z(_0307_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5083_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[3][21] ),
    .I1(\soc.spi_video_ram_1.fifo_in_address[5] ),
    .S(_2368_),
    .Z(_2372_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5084_ (.I(_2372_),
    .Z(_0308_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5085_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[3][22] ),
    .I1(\soc.spi_video_ram_1.fifo_in_address[6] ),
    .S(_2368_),
    .Z(_2373_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5086_ (.I(_2373_),
    .Z(_0309_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5087_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[3][23] ),
    .I1(\soc.spi_video_ram_1.fifo_in_address[7] ),
    .S(_2368_),
    .Z(_2374_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5088_ (.I(_2374_),
    .Z(_0310_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5089_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[3][24] ),
    .I1(\soc.spi_video_ram_1.fifo_in_address[8] ),
    .S(_2368_),
    .Z(_2375_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5090_ (.I(_2375_),
    .Z(_0311_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5091_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[3][25] ),
    .I1(\soc.spi_video_ram_1.fifo_in_address[9] ),
    .S(_2368_),
    .Z(_2376_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5092_ (.I(_2376_),
    .Z(_0312_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5093_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[3][26] ),
    .I1(\soc.spi_video_ram_1.fifo_in_address[10] ),
    .S(_2368_),
    .Z(_2377_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5094_ (.I(_2377_),
    .Z(_0313_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5095_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[3][27] ),
    .I1(\soc.spi_video_ram_1.fifo_in_address[11] ),
    .S(_2368_),
    .Z(_2378_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5096_ (.I(_2378_),
    .Z(_0314_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5097_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[3][28] ),
    .I1(\soc.spi_video_ram_1.fifo_in_address[12] ),
    .S(_2216_),
    .Z(_2379_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5098_ (.I(_2379_),
    .Z(_0315_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5099_ (.A1(_1404_),
    .A2(_1427_),
    .ZN(_2380_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5100_ (.A1(_2221_),
    .A2(_1425_),
    .ZN(_2381_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5101_ (.A1(_2380_),
    .A2(_2381_),
    .B(_1438_),
    .ZN(_2382_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5102_ (.I(\soc.rom_encoder_0.initializing_step[2] ),
    .ZN(_2383_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _5103_ (.A1(\soc.rom_encoder_0.initializing_step[4] ),
    .A2(\soc.rom_encoder_0.initializing_step[1] ),
    .A3(_1438_),
    .ZN(_2384_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5104_ (.A1(\soc.rom_encoder_0.initializing_step[3] ),
    .A2(_2383_),
    .A3(_2384_),
    .ZN(_2385_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _5105_ (.A1(_1438_),
    .A2(_2380_),
    .B(_2382_),
    .C(_2385_),
    .ZN(_2386_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5106_ (.A1(\soc.rom_encoder_0.initialized ),
    .A2(_2386_),
    .ZN(_2387_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5107_ (.A1(_0691_),
    .A2(_2387_),
    .ZN(_0316_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5108_ (.A1(_1434_),
    .A2(_1421_),
    .ZN(_2388_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _5109_ (.A1(_2223_),
    .A2(_2228_),
    .B(_2388_),
    .ZN(_2389_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5110_ (.A1(_1403_),
    .A2(_2389_),
    .ZN(_2390_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _5111_ (.A1(_1407_),
    .A2(\soc.rom_encoder_0.current_state[1] ),
    .A3(_2390_),
    .ZN(_2391_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5112_ (.I(_2391_),
    .Z(_2392_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5113_ (.I(_2391_),
    .Z(_2393_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5114_ (.I(_2225_),
    .Z(_2394_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5115_ (.I(_2394_),
    .Z(_2395_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5116_ (.A1(\soc.rom_encoder_0.request_data_out[0] ),
    .A2(_2395_),
    .ZN(_2396_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5117_ (.A1(net5),
    .A2(_2223_),
    .ZN(_2397_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5118_ (.A1(_2393_),
    .A2(_2396_),
    .A3(_2397_),
    .ZN(_2398_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5119_ (.A1(\soc.cpu.DMuxJMP.sel[0] ),
    .A2(_2392_),
    .B(_2398_),
    .ZN(_2399_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5120_ (.A1(_0691_),
    .A2(_2399_),
    .ZN(_0317_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5121_ (.I(_0690_),
    .Z(_2400_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5122_ (.A1(\soc.rom_encoder_0.request_data_out[1] ),
    .A2(_2395_),
    .ZN(_2401_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5123_ (.A1(net6),
    .A2(_2223_),
    .ZN(_2402_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5124_ (.A1(_2393_),
    .A2(_2401_),
    .A3(_2402_),
    .ZN(_2403_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5125_ (.A1(\soc.cpu.DMuxJMP.sel[1] ),
    .A2(_2392_),
    .B(_2403_),
    .ZN(_2404_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5126_ (.A1(_2400_),
    .A2(_2404_),
    .ZN(_0318_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5127_ (.A1(\soc.rom_encoder_0.request_data_out[2] ),
    .A2(_2395_),
    .ZN(_2405_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5128_ (.A1(net7),
    .A2(_2223_),
    .ZN(_2406_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5129_ (.A1(_2393_),
    .A2(_2405_),
    .A3(_2406_),
    .ZN(_2407_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5130_ (.A1(\soc.cpu.DMuxJMP.sel[2] ),
    .A2(_2392_),
    .B(_2407_),
    .ZN(_2408_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5131_ (.A1(_2400_),
    .A2(_2408_),
    .ZN(_0319_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5132_ (.A1(\soc.rom_encoder_0.request_data_out[3] ),
    .A2(_2395_),
    .ZN(_2409_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5133_ (.A1(net8),
    .A2(_2223_),
    .ZN(_2410_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5134_ (.A1(_2393_),
    .A2(_2409_),
    .A3(_2410_),
    .ZN(_2411_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5135_ (.A1(\soc.cpu.instruction[3] ),
    .A2(_2392_),
    .B(_2411_),
    .ZN(_2412_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5136_ (.A1(_2400_),
    .A2(_2412_),
    .ZN(_0320_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5137_ (.I(_2394_),
    .Z(_2413_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5138_ (.I(_2391_),
    .Z(_2414_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5139_ (.A1(\soc.rom_encoder_0.request_data_out[4] ),
    .A2(_2395_),
    .ZN(_2415_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5140_ (.A1(_2240_),
    .A2(_2413_),
    .B(_2414_),
    .C(_2415_),
    .ZN(_2416_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5141_ (.A1(\soc.cpu.instruction[4] ),
    .A2(_2392_),
    .B(_2416_),
    .ZN(_2417_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5142_ (.A1(_2400_),
    .A2(_2417_),
    .ZN(_0321_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5143_ (.A1(\soc.rom_encoder_0.request_data_out[5] ),
    .A2(_2395_),
    .ZN(_2418_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5144_ (.A1(_2245_),
    .A2(_2413_),
    .B(_2414_),
    .C(_2418_),
    .ZN(_2419_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5145_ (.A1(\soc.cpu.instruction[5] ),
    .A2(_2392_),
    .B(_2419_),
    .ZN(_2420_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5146_ (.A1(_2400_),
    .A2(_2420_),
    .ZN(_0322_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5147_ (.A1(\soc.rom_encoder_0.request_data_out[6] ),
    .A2(_2395_),
    .ZN(_2421_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5148_ (.A1(_2247_),
    .A2(_2413_),
    .B(_2414_),
    .C(_2421_),
    .ZN(_2422_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5149_ (.A1(_0990_),
    .A2(_2392_),
    .B(_2422_),
    .ZN(_2423_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5150_ (.A1(_2400_),
    .A2(_2423_),
    .ZN(_0323_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5151_ (.A1(\soc.rom_encoder_0.request_data_out[7] ),
    .A2(_2395_),
    .ZN(_2424_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5152_ (.A1(_2249_),
    .A2(_2413_),
    .B(_2414_),
    .C(_2424_),
    .ZN(_2425_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5153_ (.A1(_0954_),
    .A2(_2392_),
    .B(_2425_),
    .ZN(_2426_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5154_ (.A1(_2400_),
    .A2(_2426_),
    .ZN(_0324_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5155_ (.A1(\soc.rom_encoder_0.request_data_out[8] ),
    .A2(_2394_),
    .ZN(_2427_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5156_ (.A1(_2252_),
    .A2(_2413_),
    .B(_2414_),
    .C(_2427_),
    .ZN(_2428_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5157_ (.A1(_0926_),
    .A2(_2392_),
    .B(_2428_),
    .ZN(_2429_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5158_ (.A1(_2400_),
    .A2(_2429_),
    .ZN(_0325_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5159_ (.A1(\soc.rom_encoder_0.request_data_out[9] ),
    .A2(_2394_),
    .ZN(_2430_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5160_ (.A1(_2254_),
    .A2(_2413_),
    .B(_2414_),
    .C(_2430_),
    .ZN(_2431_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5161_ (.A1(_1011_),
    .A2(_2392_),
    .B(_2431_),
    .ZN(_2432_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5162_ (.A1(_2400_),
    .A2(_2432_),
    .ZN(_0326_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5163_ (.A1(\soc.rom_encoder_0.request_data_out[10] ),
    .A2(_2394_),
    .ZN(_2433_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5164_ (.A1(_2256_),
    .A2(_2413_),
    .B(_2414_),
    .C(_2433_),
    .ZN(_2434_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5165_ (.A1(_0923_),
    .A2(_2393_),
    .B(_2434_),
    .ZN(_2435_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5166_ (.A1(_2400_),
    .A2(_2435_),
    .ZN(_0327_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5167_ (.I(_0690_),
    .Z(_2436_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5168_ (.A1(\soc.rom_encoder_0.request_data_out[11] ),
    .A2(_2394_),
    .ZN(_2437_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5169_ (.A1(_2258_),
    .A2(_2413_),
    .B(_2414_),
    .C(_2437_),
    .ZN(_2438_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5170_ (.A1(\soc.cpu.ALU.zx ),
    .A2(_2393_),
    .B(_2438_),
    .ZN(_2439_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5171_ (.A1(_2436_),
    .A2(_2439_),
    .ZN(_0328_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5172_ (.A1(\soc.rom_encoder_0.request_data_out[12] ),
    .A2(_2394_),
    .ZN(_2440_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5173_ (.A1(_2260_),
    .A2(_2413_),
    .B(_2414_),
    .C(_2440_),
    .ZN(_2441_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5174_ (.A1(_0887_),
    .A2(_2393_),
    .B(_2441_),
    .ZN(_2442_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5175_ (.A1(_2436_),
    .A2(_2442_),
    .ZN(_0329_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5176_ (.A1(\soc.rom_encoder_0.request_data_out[13] ),
    .A2(_2394_),
    .ZN(_2443_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5177_ (.A1(_2262_),
    .A2(_2413_),
    .B(_2414_),
    .C(_2443_),
    .ZN(_2444_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5178_ (.A1(\soc.cpu.instruction[13] ),
    .A2(_2393_),
    .B(_2444_),
    .ZN(_2445_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5179_ (.A1(_2436_),
    .A2(_2445_),
    .ZN(_0330_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5180_ (.A1(\soc.rom_encoder_0.request_data_out[14] ),
    .A2(_2394_),
    .ZN(_2446_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5181_ (.A1(_2264_),
    .A2(_2395_),
    .B(_2391_),
    .C(_2446_),
    .ZN(_2447_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5182_ (.A1(\soc.cpu.instruction[14] ),
    .A2(_2393_),
    .B(_2447_),
    .ZN(_2448_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5183_ (.A1(_2436_),
    .A2(_2448_),
    .ZN(_0331_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5184_ (.A1(\soc.rom_encoder_0.request_data_out[15] ),
    .A2(_2394_),
    .ZN(_2449_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5185_ (.A1(_2266_),
    .A2(_2395_),
    .B(_2391_),
    .C(_2449_),
    .ZN(_2450_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5186_ (.A1(_0846_),
    .A2(_2393_),
    .B(_2450_),
    .ZN(_2451_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5187_ (.A1(_2436_),
    .A2(_2451_),
    .ZN(_0332_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5188_ (.A1(_1426_),
    .A2(_1408_),
    .B1(_1419_),
    .B2(_1425_),
    .ZN(_2452_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5189_ (.A1(_1410_),
    .A2(_2385_),
    .B(_2452_),
    .ZN(_2453_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5190_ (.A1(_1426_),
    .A2(_1420_),
    .ZN(_2454_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5191_ (.A1(_2390_),
    .A2(_2454_),
    .ZN(_2455_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5192_ (.I0(net62),
    .I1(_2453_),
    .S(_2455_),
    .Z(_2456_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5193_ (.A1(_1461_),
    .A2(_2456_),
    .Z(_2457_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5194_ (.I(_2457_),
    .Z(_0333_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5195_ (.A1(_1407_),
    .A2(_2224_),
    .ZN(_2458_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5196_ (.A1(_2458_),
    .A2(_2269_),
    .B(_1403_),
    .ZN(_2459_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _5197_ (.A1(_1426_),
    .A2(_2221_),
    .A3(_1424_),
    .A4(_2459_),
    .Z(_2460_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5198_ (.A1(\soc.rom_encoder_0.sram_sio_oe ),
    .A2(_2460_),
    .B(_0690_),
    .ZN(_2461_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _5199_ (.A1(_1426_),
    .A2(_1422_),
    .A3(_2459_),
    .B(_2461_),
    .ZN(_0334_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5200_ (.A1(_1412_),
    .A2(_1417_),
    .B(_2459_),
    .ZN(_2462_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5201_ (.A1(_1406_),
    .A2(_1409_),
    .A3(_2385_),
    .ZN(_2463_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5202_ (.A1(_1439_),
    .A2(_1428_),
    .ZN(_2464_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _5203_ (.A1(_2389_),
    .A2(_2462_),
    .A3(_2463_),
    .A4(_2464_),
    .ZN(_2465_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5204_ (.A1(_2230_),
    .A2(_2465_),
    .ZN(_2466_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5205_ (.A1(_1419_),
    .A2(_2466_),
    .Z(_2467_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5206_ (.A1(_2436_),
    .A2(_2467_),
    .ZN(_0335_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5207_ (.A1(_2389_),
    .A2(_2462_),
    .A3(_2463_),
    .ZN(_2468_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5208_ (.A1(_1419_),
    .A2(_2468_),
    .B(\soc.rom_encoder_0.current_state[1] ),
    .ZN(_2469_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5209_ (.A1(_1656_),
    .A2(_2465_),
    .B(_2469_),
    .C(_0676_),
    .ZN(_0336_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _5210_ (.A1(_1426_),
    .A2(_2468_),
    .B(_1428_),
    .C(_0690_),
    .ZN(_2470_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5211_ (.A1(_1413_),
    .A2(_2465_),
    .B(_2470_),
    .ZN(_0337_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5212_ (.I(_0689_),
    .Z(_2471_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _5213_ (.A1(_1438_),
    .A2(_2380_),
    .B(_2382_),
    .C(_2471_),
    .ZN(_0338_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5214_ (.A1(\soc.rom_encoder_0.initializing_step[1] ),
    .A2(_1438_),
    .ZN(_2472_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5215_ (.A1(_1410_),
    .A2(_1440_),
    .ZN(_2473_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5216_ (.A1(_2472_),
    .A2(_2473_),
    .ZN(_2474_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5217_ (.A1(_1438_),
    .A2(_2380_),
    .B(\soc.rom_encoder_0.initializing_step[1] ),
    .ZN(_2475_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _5218_ (.A1(_2380_),
    .A2(_2474_),
    .B(_2475_),
    .C(_2471_),
    .ZN(_0339_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5219_ (.A1(_1403_),
    .A2(_1409_),
    .ZN(_2476_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5220_ (.A1(\soc.rom_encoder_0.initializing_step[2] ),
    .A2(_2476_),
    .ZN(_2477_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5221_ (.A1(\soc.rom_encoder_0.initializing_step[2] ),
    .A2(\soc.rom_encoder_0.initializing_step[1] ),
    .A3(_1438_),
    .ZN(_2478_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5222_ (.A1(_1406_),
    .A2(_2380_),
    .A3(_2478_),
    .ZN(_2479_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _5223_ (.A1(_2383_),
    .A2(_2472_),
    .B1(_2477_),
    .B2(_2479_),
    .C(_0690_),
    .ZN(_0340_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5224_ (.I(\soc.rom_encoder_0.initializing_step[3] ),
    .ZN(_2480_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5225_ (.A1(\soc.rom_encoder_0.initializing_step[3] ),
    .A2(_2476_),
    .ZN(_2481_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5226_ (.A1(_2480_),
    .A2(_2478_),
    .Z(_2482_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5227_ (.A1(_1406_),
    .A2(_2380_),
    .A3(_2482_),
    .ZN(_2483_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _5228_ (.A1(_2480_),
    .A2(_2478_),
    .B1(_2481_),
    .B2(_2483_),
    .C(_0690_),
    .ZN(_0341_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5229_ (.A1(_2476_),
    .A2(_2482_),
    .ZN(_2484_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5230_ (.A1(_2221_),
    .A2(_2380_),
    .ZN(_2485_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5231_ (.A1(\soc.rom_encoder_0.initializing_step[4] ),
    .A2(_2484_),
    .B(_2485_),
    .ZN(_2486_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _5232_ (.A1(\soc.rom_encoder_0.initializing_step[4] ),
    .A2(_2484_),
    .B(_2486_),
    .C(_2471_),
    .ZN(_0342_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5233_ (.A1(_2436_),
    .A2(\soc.ram_encoder_0.toggled_sram_sck ),
    .ZN(_0343_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5234_ (.I(\soc.ram_encoder_0.input_bits_left[2] ),
    .ZN(_2487_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _5235_ (.A1(\soc.ram_encoder_0.current_state[2] ),
    .A2(_1496_),
    .Z(_2488_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _5236_ (.A1(_2487_),
    .A2(\soc.ram_encoder_0.input_bits_left[3] ),
    .A3(\soc.ram_encoder_0.input_bits_left[4] ),
    .B(_2488_),
    .ZN(_2489_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _5237_ (.A1(\soc.ram_encoder_0.current_state[2] ),
    .A2(_1490_),
    .A3(_1502_),
    .ZN(_2490_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5238_ (.A1(\soc.ram_encoder_0.request_write ),
    .A2(_1511_),
    .B(_2490_),
    .ZN(_2491_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5239_ (.A1(\soc.ram_encoder_0.toggled_sram_sck ),
    .A2(_2491_),
    .ZN(_2492_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5240_ (.A1(_1501_),
    .A2(_2489_),
    .B(_2492_),
    .ZN(_2493_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5241_ (.A1(_0674_),
    .A2(_2493_),
    .ZN(_2494_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5242_ (.A1(\soc.ram_encoder_0.input_bits_left[2] ),
    .A2(_2494_),
    .Z(_2495_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5243_ (.A1(\soc.ram_encoder_0.input_bits_left[2] ),
    .A2(_2494_),
    .ZN(_2496_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5244_ (.A1(_1489_),
    .A2(_2495_),
    .B(_2496_),
    .ZN(_0344_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5245_ (.A1(\soc.ram_encoder_0.input_bits_left[3] ),
    .A2(_2495_),
    .Z(_2497_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5246_ (.A1(_2488_),
    .A2(_2494_),
    .Z(_2498_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5247_ (.A1(\soc.ram_encoder_0.input_bits_left[3] ),
    .A2(_2495_),
    .ZN(_2499_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5248_ (.A1(_2497_),
    .A2(_2498_),
    .A3(_2499_),
    .ZN(_0345_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5249_ (.A1(\soc.ram_encoder_0.input_bits_left[4] ),
    .A2(_2497_),
    .ZN(_2500_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5250_ (.A1(\soc.ram_encoder_0.input_bits_left[4] ),
    .A2(_2497_),
    .Z(_2501_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5251_ (.A1(_2498_),
    .A2(_2500_),
    .A3(_2501_),
    .ZN(_0346_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5252_ (.I(\soc.ram_encoder_0.input_buffer[0] ),
    .ZN(_2502_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5253_ (.A1(\soc.ram_encoder_0.toggled_sram_sck ),
    .A2(_2488_),
    .ZN(_2503_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5254_ (.I(_2503_),
    .Z(_2504_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5255_ (.I(_2503_),
    .Z(_2505_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5256_ (.A1(net1),
    .A2(_2505_),
    .B(_2250_),
    .ZN(_2506_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5257_ (.A1(_2502_),
    .A2(_2504_),
    .B(_2506_),
    .ZN(_0347_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5258_ (.I(\soc.ram_encoder_0.input_buffer[1] ),
    .ZN(_2507_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5259_ (.I(_0675_),
    .Z(_2508_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5260_ (.A1(net2),
    .A2(_2505_),
    .B(_2508_),
    .ZN(_2509_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5261_ (.A1(_2507_),
    .A2(_2504_),
    .B(_2509_),
    .ZN(_0348_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5262_ (.I(\soc.ram_encoder_0.input_buffer[2] ),
    .ZN(_2510_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5263_ (.A1(net3),
    .A2(_2505_),
    .B(_2508_),
    .ZN(_2511_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5264_ (.A1(_2510_),
    .A2(_2504_),
    .B(_2511_),
    .ZN(_0349_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5265_ (.I(\soc.ram_encoder_0.input_buffer[3] ),
    .ZN(_2512_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5266_ (.A1(net4),
    .A2(_2505_),
    .B(_2508_),
    .ZN(_2513_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5267_ (.A1(_2512_),
    .A2(_2504_),
    .B(_2513_),
    .ZN(_0350_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5268_ (.I(\soc.ram_encoder_0.input_buffer[4] ),
    .ZN(_2514_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5269_ (.A1(\soc.ram_encoder_0.input_buffer[0] ),
    .A2(_2505_),
    .B(_2508_),
    .ZN(_2515_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5270_ (.A1(_2514_),
    .A2(_2504_),
    .B(_2515_),
    .ZN(_0351_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5271_ (.I(\soc.ram_encoder_0.input_buffer[5] ),
    .ZN(_2516_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5272_ (.A1(\soc.ram_encoder_0.input_buffer[1] ),
    .A2(_2505_),
    .B(_2508_),
    .ZN(_2517_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5273_ (.A1(_2516_),
    .A2(_2504_),
    .B(_2517_),
    .ZN(_0352_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5274_ (.I(\soc.ram_encoder_0.input_buffer[6] ),
    .ZN(_2518_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5275_ (.A1(\soc.ram_encoder_0.input_buffer[2] ),
    .A2(_2505_),
    .B(_2508_),
    .ZN(_2519_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5276_ (.A1(_2518_),
    .A2(_2504_),
    .B(_2519_),
    .ZN(_0353_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5277_ (.I(\soc.ram_encoder_0.input_buffer[7] ),
    .ZN(_2520_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5278_ (.A1(\soc.ram_encoder_0.input_buffer[3] ),
    .A2(_2505_),
    .B(_2508_),
    .ZN(_2521_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5279_ (.A1(_2520_),
    .A2(_2504_),
    .B(_2521_),
    .ZN(_0354_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5280_ (.I(\soc.ram_encoder_0.input_buffer[8] ),
    .ZN(_2522_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5281_ (.A1(\soc.ram_encoder_0.input_buffer[4] ),
    .A2(_2503_),
    .B(_2508_),
    .ZN(_2523_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5282_ (.A1(_2522_),
    .A2(_2504_),
    .B(_2523_),
    .ZN(_0355_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5283_ (.I(\soc.ram_encoder_0.input_buffer[9] ),
    .ZN(_2524_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5284_ (.A1(\soc.ram_encoder_0.input_buffer[5] ),
    .A2(_2503_),
    .B(_2508_),
    .ZN(_2525_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5285_ (.A1(_2524_),
    .A2(_2504_),
    .B(_2525_),
    .ZN(_0356_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5286_ (.I(\soc.ram_encoder_0.input_buffer[10] ),
    .ZN(_2526_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5287_ (.A1(\soc.ram_encoder_0.input_buffer[6] ),
    .A2(_2503_),
    .B(_2508_),
    .ZN(_2527_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5288_ (.A1(_2526_),
    .A2(_2505_),
    .B(_2527_),
    .ZN(_0357_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5289_ (.I(\soc.ram_encoder_0.input_buffer[11] ),
    .ZN(_2528_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5290_ (.A1(\soc.ram_encoder_0.input_buffer[7] ),
    .A2(_2503_),
    .B(_0675_),
    .ZN(_2529_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5291_ (.A1(_2528_),
    .A2(_2505_),
    .B(_2529_),
    .ZN(_0358_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _5292_ (.A1(_1493_),
    .A2(\soc.ram_encoder_0.current_state[1] ),
    .A3(_1488_),
    .ZN(_2530_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _5293_ (.I(_0743_),
    .ZN(_2531_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5294_ (.A1(\soc.ram_step2_read_request ),
    .A2(\soc.ram_step1_write_request ),
    .B(_2531_),
    .ZN(_2532_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5295_ (.A1(_2530_),
    .A2(_2532_),
    .ZN(_2533_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5296_ (.A1(_1493_),
    .A2(_1503_),
    .ZN(_2534_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5297_ (.A1(_1512_),
    .A2(_2533_),
    .A3(_2534_),
    .ZN(_2535_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _5298_ (.A1(_2490_),
    .A2(_2492_),
    .A3(_2535_),
    .Z(_2536_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5299_ (.I(_2536_),
    .Z(_2537_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5300_ (.I(_2537_),
    .Z(_2538_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5301_ (.A1(\soc.synch_hack_writeM ),
    .A2(_0869_),
    .ZN(_2539_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5302_ (.A1(\soc.ram_encoder_0.request_write ),
    .A2(_2538_),
    .ZN(_2540_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5303_ (.A1(_2538_),
    .A2(_2539_),
    .B(_2540_),
    .ZN(_0359_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5304_ (.I(\soc.ram_encoder_0.data_out[0] ),
    .ZN(_2541_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5305_ (.I(_2537_),
    .Z(_2542_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5306_ (.A1(\soc.ram_encoder_0.request_data_out[0] ),
    .A2(_2538_),
    .ZN(_2543_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5307_ (.A1(_2541_),
    .A2(_2542_),
    .B(_2543_),
    .ZN(_0360_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5308_ (.I(\soc.ram_encoder_0.data_out[1] ),
    .ZN(_2544_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5309_ (.I(_2537_),
    .Z(_2545_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5310_ (.A1(\soc.ram_encoder_0.request_data_out[1] ),
    .A2(_2545_),
    .ZN(_2546_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5311_ (.A1(_2544_),
    .A2(_2542_),
    .B(_2546_),
    .ZN(_0361_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5312_ (.I(\soc.ram_encoder_0.data_out[2] ),
    .ZN(_2547_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5313_ (.A1(\soc.ram_encoder_0.request_data_out[2] ),
    .A2(_2545_),
    .ZN(_2548_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5314_ (.A1(_2547_),
    .A2(_2542_),
    .B(_2548_),
    .ZN(_0362_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5315_ (.I(\soc.ram_encoder_0.data_out[3] ),
    .ZN(_2549_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5316_ (.A1(\soc.ram_encoder_0.request_data_out[3] ),
    .A2(_2545_),
    .ZN(_2550_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5317_ (.A1(_2549_),
    .A2(_2542_),
    .B(_2550_),
    .ZN(_0363_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5318_ (.I(\soc.ram_encoder_0.data_out[4] ),
    .ZN(_2551_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5319_ (.A1(\soc.ram_encoder_0.request_data_out[4] ),
    .A2(_2545_),
    .ZN(_2552_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5320_ (.A1(_2551_),
    .A2(_2542_),
    .B(_2552_),
    .ZN(_0364_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5321_ (.I(\soc.ram_encoder_0.data_out[5] ),
    .ZN(_2553_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5322_ (.A1(\soc.ram_encoder_0.request_data_out[5] ),
    .A2(_2545_),
    .ZN(_2554_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5323_ (.A1(_2553_),
    .A2(_2542_),
    .B(_2554_),
    .ZN(_0365_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5324_ (.I(\soc.ram_encoder_0.data_out[6] ),
    .ZN(_2555_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5325_ (.A1(\soc.ram_encoder_0.request_data_out[6] ),
    .A2(_2545_),
    .ZN(_2556_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5326_ (.A1(_2555_),
    .A2(_2542_),
    .B(_2556_),
    .ZN(_0366_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5327_ (.I(\soc.ram_encoder_0.data_out[7] ),
    .ZN(_2557_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5328_ (.A1(\soc.ram_encoder_0.request_data_out[7] ),
    .A2(_2545_),
    .ZN(_2558_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5329_ (.A1(_2557_),
    .A2(_2542_),
    .B(_2558_),
    .ZN(_0367_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5330_ (.I(\soc.ram_encoder_0.data_out[8] ),
    .ZN(_2559_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5331_ (.A1(\soc.ram_encoder_0.request_data_out[8] ),
    .A2(_2545_),
    .ZN(_2560_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5332_ (.A1(_2559_),
    .A2(_2542_),
    .B(_2560_),
    .ZN(_0368_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5333_ (.I(\soc.ram_encoder_0.data_out[9] ),
    .ZN(_2561_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5334_ (.A1(\soc.ram_encoder_0.request_data_out[9] ),
    .A2(_2545_),
    .ZN(_2562_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5335_ (.A1(_2561_),
    .A2(_2538_),
    .B(_2562_),
    .ZN(_0369_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5336_ (.I(\soc.ram_encoder_0.data_out[10] ),
    .ZN(_2563_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5337_ (.A1(\soc.ram_encoder_0.request_data_out[10] ),
    .A2(_2545_),
    .ZN(_2564_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5338_ (.A1(_2563_),
    .A2(_2538_),
    .B(_2564_),
    .ZN(_0370_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5339_ (.I(\soc.ram_encoder_0.data_out[11] ),
    .ZN(_2565_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 _5340_ (.I(_2537_),
    .Z(_2566_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5341_ (.A1(\soc.ram_encoder_0.request_data_out[11] ),
    .A2(_2566_),
    .ZN(_2567_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5342_ (.A1(_2565_),
    .A2(_2538_),
    .B(_2567_),
    .ZN(_0371_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5343_ (.I(\soc.ram_encoder_0.data_out[12] ),
    .ZN(_2568_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5344_ (.A1(\soc.ram_encoder_0.request_data_out[12] ),
    .A2(_2566_),
    .ZN(_2569_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5345_ (.A1(_2568_),
    .A2(_2538_),
    .B(_2569_),
    .ZN(_0372_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5346_ (.I(\soc.ram_encoder_0.data_out[13] ),
    .ZN(_2570_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5347_ (.A1(\soc.ram_encoder_0.request_data_out[13] ),
    .A2(_2566_),
    .ZN(_2571_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5348_ (.A1(_2570_),
    .A2(_2538_),
    .B(_2571_),
    .ZN(_0373_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5349_ (.I(\soc.ram_encoder_0.data_out[14] ),
    .ZN(_2572_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5350_ (.A1(\soc.ram_encoder_0.request_data_out[14] ),
    .A2(_2566_),
    .ZN(_2573_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5351_ (.A1(_2572_),
    .A2(_2538_),
    .B(_2573_),
    .ZN(_0374_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5352_ (.I(\soc.ram_encoder_0.data_out[15] ),
    .ZN(_2574_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5353_ (.A1(\soc.ram_encoder_0.request_data_out[15] ),
    .A2(_2566_),
    .ZN(_2575_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5354_ (.A1(_2574_),
    .A2(_2538_),
    .B(_2575_),
    .ZN(_0375_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5355_ (.I0(\soc.ram_encoder_0.address[0] ),
    .I1(\soc.ram_encoder_0.request_address[0] ),
    .S(_2566_),
    .Z(_2576_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5356_ (.I(_2576_),
    .Z(_0376_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5357_ (.I0(\soc.ram_encoder_0.address[1] ),
    .I1(\soc.ram_encoder_0.request_address[1] ),
    .S(_2566_),
    .Z(_2577_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5358_ (.I(_2577_),
    .Z(_0377_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5359_ (.I0(\soc.ram_encoder_0.address[2] ),
    .I1(\soc.ram_encoder_0.request_address[2] ),
    .S(_2566_),
    .Z(_2578_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5360_ (.I(_2578_),
    .Z(_0378_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5361_ (.I0(\soc.ram_encoder_0.address[3] ),
    .I1(\soc.ram_encoder_0.request_address[3] ),
    .S(_2566_),
    .Z(_2579_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5362_ (.I(_2579_),
    .Z(_0379_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5363_ (.I0(\soc.ram_encoder_0.address[4] ),
    .I1(\soc.ram_encoder_0.request_address[4] ),
    .S(_2566_),
    .Z(_2580_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5364_ (.I(_2580_),
    .Z(_0380_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _5365_ (.I(_2537_),
    .Z(_2581_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5366_ (.I0(\soc.ram_encoder_0.address[5] ),
    .I1(\soc.ram_encoder_0.request_address[5] ),
    .S(_2581_),
    .Z(_2582_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5367_ (.I(_2582_),
    .Z(_0381_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5368_ (.I0(\soc.ram_encoder_0.address[6] ),
    .I1(\soc.ram_encoder_0.request_address[6] ),
    .S(_2581_),
    .Z(_2583_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5369_ (.I(_2583_),
    .Z(_0382_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5370_ (.I0(\soc.ram_encoder_0.address[7] ),
    .I1(\soc.ram_encoder_0.request_address[7] ),
    .S(_2581_),
    .Z(_2584_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5371_ (.I(_2584_),
    .Z(_0383_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5372_ (.I0(\soc.ram_encoder_0.address[8] ),
    .I1(\soc.ram_encoder_0.request_address[8] ),
    .S(_2581_),
    .Z(_2585_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5373_ (.I(_2585_),
    .Z(_0384_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5374_ (.I0(\soc.ram_encoder_0.address[9] ),
    .I1(\soc.ram_encoder_0.request_address[9] ),
    .S(_2581_),
    .Z(_2586_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5375_ (.I(_2586_),
    .Z(_0385_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5376_ (.I0(\soc.ram_encoder_0.address[10] ),
    .I1(\soc.ram_encoder_0.request_address[10] ),
    .S(_2581_),
    .Z(_2587_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5377_ (.I(_2587_),
    .Z(_0386_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5378_ (.I0(\soc.ram_encoder_0.address[11] ),
    .I1(\soc.ram_encoder_0.request_address[11] ),
    .S(_2581_),
    .Z(_2588_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5379_ (.I(_2588_),
    .Z(_0387_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5380_ (.I0(\soc.ram_encoder_0.address[12] ),
    .I1(\soc.ram_encoder_0.request_address[12] ),
    .S(_2581_),
    .Z(_2589_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5381_ (.I(_2589_),
    .Z(_0388_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5382_ (.I0(\soc.ram_encoder_0.address[13] ),
    .I1(\soc.ram_encoder_0.request_address[13] ),
    .S(_2581_),
    .Z(_2590_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5383_ (.I(_2590_),
    .Z(_0389_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5384_ (.I0(\soc.ram_encoder_0.address[14] ),
    .I1(\soc.ram_encoder_0.request_address[14] ),
    .S(_2581_),
    .Z(_2591_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5385_ (.I(_2591_),
    .Z(_0390_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5386_ (.A1(\soc.ram_encoder_0.initializing_step[4] ),
    .A2(\soc.ram_encoder_0.initializing_step[2] ),
    .ZN(_2592_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5387_ (.A1(\soc.ram_encoder_0.initializing_step[1] ),
    .A2(\soc.ram_encoder_0.initializing_step[0] ),
    .ZN(_2593_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5388_ (.A1(\soc.ram_encoder_0.initializing_step[3] ),
    .A2(_2592_),
    .A3(_2593_),
    .ZN(_2594_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5389_ (.A1(\soc.ram_encoder_0.toggled_sram_sck ),
    .A2(_1491_),
    .ZN(_2595_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5390_ (.A1(_1495_),
    .A2(_2595_),
    .ZN(_2596_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5391_ (.A1(_1405_),
    .A2(_2334_),
    .ZN(_2597_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5392_ (.A1(\soc.ram_encoder_0.initializing_step[0] ),
    .A2(_2597_),
    .ZN(_2598_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5393_ (.A1(\soc.ram_encoder_0.initializing_step[0] ),
    .A2(_2596_),
    .B(_2598_),
    .ZN(_2599_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5394_ (.A1(\soc.ram_encoder_0.initialized ),
    .A2(_1955_),
    .ZN(_2600_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _5395_ (.A1(_1461_),
    .A2(_2594_),
    .A3(_2599_),
    .B(_2600_),
    .ZN(_0391_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _5396_ (.A1(_1504_),
    .A2(_1499_),
    .B(_2489_),
    .C(\soc.ram_encoder_0.toggled_sram_sck ),
    .ZN(_2601_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _5397_ (.A1(_1489_),
    .A2(\soc.ram_encoder_0.current_state[1] ),
    .A3(_2601_),
    .ZN(_2602_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5398_ (.I(_2602_),
    .Z(_2603_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5399_ (.I(_2602_),
    .Z(_2604_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5400_ (.A1(_1493_),
    .A2(_1496_),
    .ZN(_2605_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5401_ (.I(_2605_),
    .Z(_2606_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5402_ (.A1(\soc.ram_encoder_0.request_data_out[0] ),
    .A2(_2606_),
    .ZN(_2607_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5403_ (.A1(net1),
    .A2(_2488_),
    .ZN(_2608_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5404_ (.A1(_2604_),
    .A2(_2607_),
    .A3(_2608_),
    .ZN(_2609_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5405_ (.A1(\soc.ram_data_out[0] ),
    .A2(_2603_),
    .B(_2609_),
    .ZN(_2610_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5406_ (.A1(_2436_),
    .A2(_2610_),
    .ZN(_0392_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5407_ (.A1(\soc.ram_encoder_0.request_data_out[1] ),
    .A2(_2606_),
    .ZN(_2611_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5408_ (.A1(net2),
    .A2(_2488_),
    .ZN(_2612_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5409_ (.A1(_2604_),
    .A2(_2611_),
    .A3(_2612_),
    .ZN(_2613_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5410_ (.A1(\soc.ram_data_out[1] ),
    .A2(_2603_),
    .B(_2613_),
    .ZN(_2614_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5411_ (.A1(_2436_),
    .A2(_2614_),
    .ZN(_0393_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5412_ (.I(_0689_),
    .Z(_2615_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5413_ (.A1(\soc.ram_encoder_0.request_data_out[2] ),
    .A2(_2606_),
    .ZN(_2616_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5414_ (.A1(net3),
    .A2(_2488_),
    .ZN(_2617_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5415_ (.A1(_2604_),
    .A2(_2616_),
    .A3(_2617_),
    .ZN(_2618_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5416_ (.A1(\soc.ram_data_out[2] ),
    .A2(_2603_),
    .B(_2618_),
    .ZN(_2619_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5417_ (.A1(_2615_),
    .A2(_2619_),
    .ZN(_0394_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5418_ (.A1(\soc.ram_encoder_0.request_data_out[3] ),
    .A2(_2606_),
    .ZN(_2620_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5419_ (.A1(net4),
    .A2(_2488_),
    .ZN(_2621_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5420_ (.A1(_2604_),
    .A2(_2620_),
    .A3(_2621_),
    .ZN(_2622_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5421_ (.A1(\soc.ram_data_out[3] ),
    .A2(_2603_),
    .B(_2622_),
    .ZN(_2623_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5422_ (.A1(_2615_),
    .A2(_2623_),
    .ZN(_0395_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5423_ (.I(_2605_),
    .Z(_2624_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5424_ (.I(_2602_),
    .Z(_2625_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5425_ (.A1(\soc.ram_encoder_0.request_data_out[4] ),
    .A2(_2606_),
    .ZN(_2626_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5426_ (.A1(_2502_),
    .A2(_2624_),
    .B(_2625_),
    .C(_2626_),
    .ZN(_2627_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5427_ (.A1(\soc.ram_data_out[4] ),
    .A2(_2603_),
    .B(_2627_),
    .ZN(_2628_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5428_ (.A1(_2615_),
    .A2(_2628_),
    .ZN(_0396_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5429_ (.A1(\soc.ram_encoder_0.request_data_out[5] ),
    .A2(_2606_),
    .ZN(_2629_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5430_ (.A1(_2507_),
    .A2(_2624_),
    .B(_2625_),
    .C(_2629_),
    .ZN(_2630_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5431_ (.A1(\soc.ram_data_out[5] ),
    .A2(_2603_),
    .B(_2630_),
    .ZN(_2631_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5432_ (.A1(_2615_),
    .A2(_2631_),
    .ZN(_0397_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5433_ (.A1(\soc.ram_encoder_0.request_data_out[6] ),
    .A2(_2606_),
    .ZN(_2632_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5434_ (.A1(_2510_),
    .A2(_2624_),
    .B(_2625_),
    .C(_2632_),
    .ZN(_2633_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5435_ (.A1(\soc.ram_data_out[6] ),
    .A2(_2603_),
    .B(_2633_),
    .ZN(_2634_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5436_ (.A1(_2615_),
    .A2(_2634_),
    .ZN(_0398_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5437_ (.A1(\soc.ram_encoder_0.request_data_out[7] ),
    .A2(_2606_),
    .ZN(_2635_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5438_ (.A1(_2512_),
    .A2(_2624_),
    .B(_2625_),
    .C(_2635_),
    .ZN(_2636_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5439_ (.A1(\soc.ram_data_out[7] ),
    .A2(_2603_),
    .B(_2636_),
    .ZN(_2637_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5440_ (.A1(_2615_),
    .A2(_2637_),
    .ZN(_0399_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5441_ (.A1(\soc.ram_encoder_0.request_data_out[8] ),
    .A2(_2605_),
    .ZN(_2638_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5442_ (.A1(_2514_),
    .A2(_2624_),
    .B(_2625_),
    .C(_2638_),
    .ZN(_2639_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5443_ (.A1(\soc.ram_data_out[8] ),
    .A2(_2603_),
    .B(_2639_),
    .ZN(_2640_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5444_ (.A1(_2615_),
    .A2(_2640_),
    .ZN(_0400_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5445_ (.A1(\soc.ram_encoder_0.request_data_out[9] ),
    .A2(_2605_),
    .ZN(_2641_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5446_ (.A1(_2516_),
    .A2(_2624_),
    .B(_2625_),
    .C(_2641_),
    .ZN(_2642_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5447_ (.A1(\soc.ram_data_out[9] ),
    .A2(_2603_),
    .B(_2642_),
    .ZN(_2643_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5448_ (.A1(_2615_),
    .A2(_2643_),
    .ZN(_0401_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5449_ (.A1(\soc.ram_encoder_0.request_data_out[10] ),
    .A2(_2605_),
    .ZN(_2644_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5450_ (.A1(_2518_),
    .A2(_2624_),
    .B(_2625_),
    .C(_2644_),
    .ZN(_2645_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5451_ (.A1(\soc.ram_data_out[10] ),
    .A2(_2604_),
    .B(_2645_),
    .ZN(_2646_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5452_ (.A1(_2615_),
    .A2(_2646_),
    .ZN(_0402_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5453_ (.A1(\soc.ram_encoder_0.request_data_out[11] ),
    .A2(_2605_),
    .ZN(_2647_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5454_ (.A1(_2520_),
    .A2(_2624_),
    .B(_2625_),
    .C(_2647_),
    .ZN(_2648_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5455_ (.A1(\soc.ram_data_out[11] ),
    .A2(_2604_),
    .B(_2648_),
    .ZN(_2649_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5456_ (.A1(_2615_),
    .A2(_2649_),
    .ZN(_0403_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5457_ (.A1(\soc.ram_encoder_0.request_data_out[12] ),
    .A2(_2605_),
    .ZN(_2650_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5458_ (.A1(_2522_),
    .A2(_2624_),
    .B(_2625_),
    .C(_2650_),
    .ZN(_2651_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5459_ (.A1(\soc.ram_data_out[12] ),
    .A2(_2604_),
    .B(_2651_),
    .ZN(_2652_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5460_ (.A1(_2471_),
    .A2(_2652_),
    .ZN(_0404_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5461_ (.A1(\soc.ram_encoder_0.request_data_out[13] ),
    .A2(_2605_),
    .ZN(_2653_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5462_ (.A1(_2524_),
    .A2(_2624_),
    .B(_2625_),
    .C(_2653_),
    .ZN(_2654_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5463_ (.A1(\soc.ram_data_out[13] ),
    .A2(_2604_),
    .B(_2654_),
    .ZN(_2655_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5464_ (.A1(_2471_),
    .A2(_2655_),
    .ZN(_0405_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5465_ (.A1(\soc.ram_encoder_0.request_data_out[14] ),
    .A2(_2605_),
    .ZN(_2656_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5466_ (.A1(_2526_),
    .A2(_2606_),
    .B(_2602_),
    .C(_2656_),
    .ZN(_2657_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5467_ (.A1(\soc.ram_data_out[14] ),
    .A2(_2604_),
    .B(_2657_),
    .ZN(_2658_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5468_ (.A1(_2471_),
    .A2(_2658_),
    .ZN(_0406_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5469_ (.A1(\soc.ram_encoder_0.request_data_out[15] ),
    .A2(_2605_),
    .ZN(_2659_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5470_ (.A1(_2528_),
    .A2(_2606_),
    .B(_2602_),
    .C(_2659_),
    .ZN(_2660_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5471_ (.A1(\soc.ram_data_out[15] ),
    .A2(_2604_),
    .B(_2660_),
    .ZN(_2661_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5472_ (.A1(_2471_),
    .A2(_2661_),
    .ZN(_0407_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5473_ (.A1(_2534_),
    .A2(_2601_),
    .Z(_2662_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5474_ (.A1(_1492_),
    .A2(_2594_),
    .ZN(_2663_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _5475_ (.A1(_1493_),
    .A2(_1490_),
    .B(_1495_),
    .C(_2663_),
    .ZN(_2664_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5476_ (.A1(net81),
    .A2(_2662_),
    .B(_0690_),
    .ZN(_2665_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5477_ (.A1(_2662_),
    .A2(_2664_),
    .B(_2665_),
    .ZN(_0408_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5478_ (.A1(_2492_),
    .A2(_2535_),
    .B(\soc.ram_encoder_0.sram_sio_oe ),
    .ZN(_2666_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5479_ (.A1(_1955_),
    .A2(_2542_),
    .A3(_2666_),
    .ZN(_0409_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5480_ (.A1(_1502_),
    .A2(_2594_),
    .ZN(_2667_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _5481_ (.A1(_2334_),
    .A2(_1495_),
    .A3(_2667_),
    .ZN(_2668_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5482_ (.A1(_1517_),
    .A2(_2533_),
    .ZN(_2669_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _5483_ (.A1(_2601_),
    .A2(_2668_),
    .A3(_2669_),
    .ZN(_2670_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5484_ (.A1(_1512_),
    .A2(_2670_),
    .ZN(_2671_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _5485_ (.A1(\soc.ram_encoder_0.request_write ),
    .A2(_2490_),
    .B(_2530_),
    .C(_2671_),
    .ZN(_2672_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5486_ (.A1(_1488_),
    .A2(_2670_),
    .B(_1955_),
    .ZN(_2673_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5487_ (.A1(_2672_),
    .A2(_2673_),
    .ZN(_0410_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5488_ (.A1(\soc.ram_encoder_0.current_state[1] ),
    .A2(_2670_),
    .B1(_2671_),
    .B2(_1557_),
    .ZN(_2674_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5489_ (.A1(_0676_),
    .A2(_2674_),
    .ZN(_0411_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _5490_ (.A1(_2490_),
    .A2(_2670_),
    .B1(_2671_),
    .B2(_1493_),
    .C(_0690_),
    .ZN(_2675_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5491_ (.I(_2675_),
    .ZN(_0412_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5492_ (.A1(_2436_),
    .A2(_2599_),
    .ZN(_0413_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5493_ (.A1(_1488_),
    .A2(_2595_),
    .ZN(_2676_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5494_ (.A1(\soc.ram_encoder_0.initializing_step[1] ),
    .A2(_2598_),
    .Z(_2677_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _5495_ (.A1(_1516_),
    .A2(_2676_),
    .B(_2677_),
    .C(_2471_),
    .ZN(_0414_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _5496_ (.A1(\soc.ram_encoder_0.initializing_step[1] ),
    .A2(\soc.ram_encoder_0.initializing_step[0] ),
    .A3(_2597_),
    .Z(_2678_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _5497_ (.A1(_1488_),
    .A2(_2595_),
    .B1(_2678_),
    .B2(\soc.ram_encoder_0.initializing_step[2] ),
    .C(_0675_),
    .ZN(_2679_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5498_ (.A1(\soc.ram_encoder_0.initializing_step[2] ),
    .A2(_2678_),
    .B(_2679_),
    .ZN(_0415_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5499_ (.A1(\soc.ram_encoder_0.initializing_step[3] ),
    .A2(\soc.ram_encoder_0.initializing_step[2] ),
    .A3(_2678_),
    .ZN(_2680_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5500_ (.A1(_1488_),
    .A2(_2595_),
    .B(_0675_),
    .ZN(_2681_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5501_ (.A1(\soc.ram_encoder_0.initializing_step[2] ),
    .A2(_2678_),
    .B(\soc.ram_encoder_0.initializing_step[3] ),
    .ZN(_2682_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5502_ (.A1(_2681_),
    .A2(_2682_),
    .ZN(_2683_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5503_ (.A1(_2680_),
    .A2(_2683_),
    .Z(_2684_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5504_ (.I(_2684_),
    .Z(_0416_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5505_ (.A1(\soc.ram_encoder_0.initializing_step[4] ),
    .A2(_2680_),
    .Z(_2685_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5506_ (.A1(_2681_),
    .A2(_2685_),
    .ZN(_0417_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5507_ (.I(\soc.hack_clock_0.counter[0] ),
    .ZN(_2686_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5508_ (.I(\soc.hack_clock_0.counter[5] ),
    .ZN(_2687_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _5509_ (.A1(\soc.hack_clock_0.counter[4] ),
    .A2(_2687_),
    .A3(\soc.hack_clock_0.counter[6] ),
    .ZN(_2688_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5510_ (.A1(\soc.hack_clock_0.counter[3] ),
    .A2(\soc.hack_clock_0.counter[2] ),
    .ZN(_2689_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _5511_ (.A1(_2686_),
    .A2(\soc.hack_clock_0.counter[1] ),
    .A3(_2688_),
    .A4(_2689_),
    .ZN(_2690_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5512_ (.A1(_0675_),
    .A2(_2690_),
    .ZN(_2691_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5513_ (.A1(\soc.hack_clock_0.counter[0] ),
    .A2(_2691_),
    .ZN(_0418_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5514_ (.A1(\soc.hack_clock_0.counter[0] ),
    .A2(\soc.hack_clock_0.counter[1] ),
    .ZN(_2692_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5515_ (.A1(\soc.hack_clock_0.counter[0] ),
    .A2(\soc.hack_clock_0.counter[1] ),
    .Z(_2693_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _5516_ (.A1(_2691_),
    .A2(_2692_),
    .A3(_2693_),
    .ZN(_0419_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5517_ (.A1(\soc.hack_clock_0.counter[2] ),
    .A2(_2693_),
    .Z(_2694_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5518_ (.A1(\soc.hack_clock_0.counter[2] ),
    .A2(_2693_),
    .ZN(_2695_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _5519_ (.A1(_2691_),
    .A2(_2694_),
    .A3(_2695_),
    .ZN(_0420_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5520_ (.A1(\soc.hack_clock_0.counter[3] ),
    .A2(_2694_),
    .Z(_2696_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5521_ (.A1(\soc.hack_clock_0.counter[3] ),
    .A2(_2694_),
    .ZN(_2697_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _5522_ (.A1(_2691_),
    .A2(_2696_),
    .A3(_2697_),
    .ZN(_0421_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5523_ (.A1(\soc.hack_clock_0.counter[4] ),
    .A2(_2696_),
    .Z(_2698_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5524_ (.A1(\soc.hack_clock_0.counter[4] ),
    .A2(_2696_),
    .ZN(_2699_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _5525_ (.A1(_2691_),
    .A2(_2698_),
    .A3(_2699_),
    .ZN(_0422_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5526_ (.A1(_2687_),
    .A2(_2698_),
    .Z(_2700_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5527_ (.A1(_2691_),
    .A2(_2700_),
    .ZN(_0423_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5528_ (.A1(\soc.hack_clock_0.counter[5] ),
    .A2(_2698_),
    .ZN(_2701_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5529_ (.A1(\soc.hack_clock_0.counter[6] ),
    .A2(_2701_),
    .Z(_2702_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5530_ (.A1(_2691_),
    .A2(_2702_),
    .ZN(_0424_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _5531_ (.I(_0694_),
    .ZN(_2703_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _5532_ (.A1(\soc.spi_video_ram_1.write_fifo.write_pointer[2] ),
    .A2(_2703_),
    .A3(_0698_),
    .ZN(_2704_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 _5533_ (.I(_2704_),
    .Z(_2705_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5534_ (.I0(\soc.spi_video_ram_1.fifo_in_data[0] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[5][0] ),
    .S(_2705_),
    .Z(_2706_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5535_ (.I(_2706_),
    .Z(_0425_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5536_ (.I(_2704_),
    .Z(_2707_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5537_ (.I(_2704_),
    .Z(_2708_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5538_ (.A1(\soc.spi_video_ram_1.fifo_in_data[1] ),
    .A2(_2708_),
    .ZN(_2709_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5539_ (.A1(_1705_),
    .A2(_2707_),
    .B(_2709_),
    .ZN(_0426_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5540_ (.I0(\soc.spi_video_ram_1.fifo_in_data[2] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[5][2] ),
    .S(_2705_),
    .Z(_2710_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5541_ (.I(_2710_),
    .Z(_0427_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5542_ (.I0(\soc.spi_video_ram_1.fifo_in_data[3] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[5][3] ),
    .S(_2705_),
    .Z(_2711_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5543_ (.I(_2711_),
    .Z(_0428_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5544_ (.I0(\soc.spi_video_ram_1.fifo_in_data[4] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[5][4] ),
    .S(_2705_),
    .Z(_2712_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5545_ (.I(_2712_),
    .Z(_0429_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5546_ (.A1(\soc.spi_video_ram_1.fifo_in_data[5] ),
    .A2(_2708_),
    .ZN(_2713_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5547_ (.A1(_1740_),
    .A2(_2707_),
    .B(_2713_),
    .ZN(_0430_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5548_ (.I0(\soc.spi_video_ram_1.fifo_in_data[6] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[5][6] ),
    .S(_2705_),
    .Z(_2714_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5549_ (.I(_2714_),
    .Z(_0431_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5550_ (.A1(\soc.spi_video_ram_1.fifo_in_data[7] ),
    .A2(_2708_),
    .ZN(_2715_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5551_ (.A1(_1767_),
    .A2(_2707_),
    .B(_2715_),
    .ZN(_0432_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5552_ (.A1(\soc.spi_video_ram_1.fifo_in_data[8] ),
    .A2(_2708_),
    .ZN(_2716_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5553_ (.A1(_1787_),
    .A2(_2707_),
    .B(_2716_),
    .ZN(_0433_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5554_ (.A1(\soc.spi_video_ram_1.fifo_in_data[9] ),
    .A2(_2708_),
    .ZN(_2717_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5555_ (.A1(_1804_),
    .A2(_2707_),
    .B(_2717_),
    .ZN(_0434_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5556_ (.I0(\soc.spi_video_ram_1.fifo_in_data[10] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[5][10] ),
    .S(_2705_),
    .Z(_2718_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5557_ (.I(_2718_),
    .Z(_0435_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _5558_ (.I(_2704_),
    .Z(_2719_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5559_ (.I0(\soc.spi_video_ram_1.fifo_in_data[11] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[5][11] ),
    .S(_2719_),
    .Z(_2720_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5560_ (.I(_2720_),
    .Z(_0436_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5561_ (.I0(\soc.spi_video_ram_1.fifo_in_data[12] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[5][12] ),
    .S(_2719_),
    .Z(_2721_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5562_ (.I(_2721_),
    .Z(_0437_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5563_ (.A1(\soc.spi_video_ram_1.fifo_in_data[13] ),
    .A2(_2708_),
    .ZN(_2722_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5564_ (.A1(_1866_),
    .A2(_2707_),
    .B(_2722_),
    .ZN(_0438_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5565_ (.A1(\soc.spi_video_ram_1.fifo_in_data[14] ),
    .A2(_2708_),
    .ZN(_2723_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5566_ (.A1(_1889_),
    .A2(_2707_),
    .B(_2723_),
    .ZN(_0439_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5567_ (.I0(\soc.spi_video_ram_1.fifo_in_data[15] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[5][15] ),
    .S(_2719_),
    .Z(_2724_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5568_ (.I(_2724_),
    .Z(_0440_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5569_ (.A1(\soc.spi_video_ram_1.fifo_in_address[0] ),
    .A2(_2708_),
    .ZN(_2725_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5570_ (.A1(_1597_),
    .A2(_2707_),
    .B(_2725_),
    .ZN(_0441_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5571_ (.A1(\soc.spi_video_ram_1.fifo_in_address[1] ),
    .A2(_2705_),
    .ZN(_2726_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5572_ (.A1(_1625_),
    .A2(_2707_),
    .B(_2726_),
    .ZN(_0442_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5573_ (.A1(\soc.spi_video_ram_1.fifo_in_address[2] ),
    .A2(_2705_),
    .ZN(_2727_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5574_ (.A1(_1615_),
    .A2(_2707_),
    .B(_2727_),
    .ZN(_0443_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5575_ (.A1(\soc.spi_video_ram_1.fifo_in_address[3] ),
    .A2(_2705_),
    .ZN(_2728_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5576_ (.A1(_1940_),
    .A2(_2708_),
    .B(_2728_),
    .ZN(_0444_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5577_ (.A1(\soc.spi_video_ram_1.fifo_in_address[4] ),
    .A2(_2705_),
    .ZN(_2729_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5578_ (.A1(_1930_),
    .A2(_2708_),
    .B(_2729_),
    .ZN(_0445_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5579_ (.I0(\soc.spi_video_ram_1.fifo_in_address[5] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[5][21] ),
    .S(_2719_),
    .Z(_2730_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5580_ (.I(_2730_),
    .Z(_0446_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5581_ (.I0(\soc.spi_video_ram_1.fifo_in_address[6] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[5][22] ),
    .S(_2719_),
    .Z(_2731_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5582_ (.I(_2731_),
    .Z(_0447_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5583_ (.I0(\soc.spi_video_ram_1.fifo_in_address[7] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[5][23] ),
    .S(_2719_),
    .Z(_2732_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5584_ (.I(_2732_),
    .Z(_0448_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5585_ (.I0(\soc.spi_video_ram_1.fifo_in_address[8] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[5][24] ),
    .S(_2719_),
    .Z(_2733_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5586_ (.I(_2733_),
    .Z(_0449_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5587_ (.I0(\soc.spi_video_ram_1.fifo_in_address[9] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[5][25] ),
    .S(_2719_),
    .Z(_2734_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5588_ (.I(_2734_),
    .Z(_0450_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5589_ (.I0(\soc.spi_video_ram_1.fifo_in_address[10] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[5][26] ),
    .S(_2719_),
    .Z(_2735_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5590_ (.I(_2735_),
    .Z(_0451_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5591_ (.I0(\soc.spi_video_ram_1.fifo_in_address[11] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[5][27] ),
    .S(_2719_),
    .Z(_2736_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5592_ (.I(_2736_),
    .Z(_0452_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5593_ (.I0(\soc.spi_video_ram_1.fifo_in_address[12] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[5][28] ),
    .S(_2704_),
    .Z(_2737_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5594_ (.I(_2737_),
    .Z(_0453_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5595_ (.A1(\soc.rom_encoder_0.initialized ),
    .A2(_2268_),
    .ZN(_2738_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5596_ (.A1(\soc.rom_encoder_0.write_enable ),
    .A2(net45),
    .ZN(_2739_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _5597_ (.A1(\soc.rom_loader.wait_fall_clk ),
    .A2(\soc.rom_loader.writing ),
    .A3(_2738_),
    .A4(_2739_),
    .ZN(_2740_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5598_ (.A1(\soc.rom_loader.rom_request ),
    .A2(_2740_),
    .B(_2268_),
    .ZN(_2741_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5599_ (.A1(_2471_),
    .A2(_2741_),
    .ZN(_0454_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5600_ (.A1(\soc.rom_loader.rom_request ),
    .A2(_2458_),
    .B(\soc.rom_loader.writing ),
    .ZN(_2742_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _5601_ (.A1(\soc.rom_loader.writing ),
    .A2(\soc.rom_loader.was_loading ),
    .A3(_2268_),
    .Z(_2743_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5602_ (.I(_2743_),
    .Z(_0473_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _5603_ (.A1(_1461_),
    .A2(_2742_),
    .A3(_0473_),
    .ZN(_0455_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5604_ (.A1(_1403_),
    .A2(_0691_),
    .ZN(_0456_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5605_ (.A1(\soc.rom_loader.current_address[0] ),
    .A2(_0473_),
    .Z(_2744_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5606_ (.A1(_2089_),
    .A2(\soc.rom_loader.was_loading ),
    .ZN(_2745_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5607_ (.I(_2745_),
    .Z(_2746_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5608_ (.A1(\soc.rom_loader.current_address[0] ),
    .A2(_0473_),
    .ZN(_2747_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _5609_ (.A1(_2744_),
    .A2(_2746_),
    .A3(_2747_),
    .ZN(_0457_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5610_ (.A1(\soc.rom_loader.current_address[1] ),
    .A2(_2744_),
    .B(_2745_),
    .ZN(_2748_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5611_ (.A1(\soc.rom_loader.current_address[1] ),
    .A2(_2744_),
    .B(_2748_),
    .ZN(_2749_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5612_ (.I(_2749_),
    .ZN(_0458_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5613_ (.A1(\soc.rom_loader.current_address[1] ),
    .A2(_2744_),
    .B(\soc.rom_loader.current_address[2] ),
    .ZN(_2750_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _5614_ (.A1(\soc.rom_loader.current_address[2] ),
    .A2(\soc.rom_loader.current_address[1] ),
    .A3(_2744_),
    .Z(_2751_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _5615_ (.A1(_2746_),
    .A2(_2750_),
    .A3(_2751_),
    .ZN(_0459_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5616_ (.A1(\soc.rom_loader.current_address[3] ),
    .A2(_2751_),
    .ZN(_2752_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5617_ (.A1(\soc.rom_loader.current_address[3] ),
    .A2(_2751_),
    .Z(_2753_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _5618_ (.A1(_2746_),
    .A2(_2752_),
    .A3(_2753_),
    .ZN(_0460_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5619_ (.A1(\soc.rom_loader.current_address[4] ),
    .A2(_2753_),
    .ZN(_2754_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5620_ (.A1(\soc.rom_loader.current_address[4] ),
    .A2(_2753_),
    .Z(_2755_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _5621_ (.A1(_2746_),
    .A2(_2754_),
    .A3(_2755_),
    .ZN(_0461_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5622_ (.A1(\soc.rom_loader.current_address[5] ),
    .A2(_2755_),
    .ZN(_2756_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5623_ (.A1(\soc.rom_loader.current_address[5] ),
    .A2(_2755_),
    .Z(_2757_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _5624_ (.A1(_2746_),
    .A2(_2756_),
    .A3(_2757_),
    .ZN(_0462_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5625_ (.A1(\soc.rom_loader.current_address[6] ),
    .A2(_2757_),
    .ZN(_2758_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5626_ (.A1(\soc.rom_loader.current_address[6] ),
    .A2(_2757_),
    .Z(_2759_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _5627_ (.A1(_2746_),
    .A2(_2758_),
    .A3(_2759_),
    .ZN(_0463_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5628_ (.A1(\soc.rom_loader.current_address[7] ),
    .A2(_2759_),
    .B(_2745_),
    .ZN(_2760_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5629_ (.A1(\soc.rom_loader.current_address[7] ),
    .A2(_2759_),
    .B(_2760_),
    .ZN(_2761_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5630_ (.I(_2761_),
    .ZN(_0464_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5631_ (.A1(\soc.rom_loader.current_address[7] ),
    .A2(_2759_),
    .B(\soc.rom_loader.current_address[8] ),
    .ZN(_2762_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _5632_ (.A1(\soc.rom_loader.current_address[8] ),
    .A2(\soc.rom_loader.current_address[7] ),
    .A3(_2759_),
    .Z(_2763_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _5633_ (.A1(_2746_),
    .A2(_2762_),
    .A3(_2763_),
    .ZN(_0465_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5634_ (.A1(\soc.rom_loader.current_address[9] ),
    .A2(_2763_),
    .ZN(_2764_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5635_ (.A1(\soc.rom_loader.current_address[9] ),
    .A2(_2763_),
    .Z(_2765_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _5636_ (.A1(_2746_),
    .A2(_2764_),
    .A3(_2765_),
    .ZN(_0466_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5637_ (.A1(\soc.rom_loader.current_address[10] ),
    .A2(_2765_),
    .ZN(_2766_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5638_ (.A1(\soc.rom_loader.current_address[10] ),
    .A2(_2765_),
    .Z(_2767_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _5639_ (.A1(_2746_),
    .A2(_2766_),
    .A3(_2767_),
    .ZN(_0467_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5640_ (.A1(\soc.rom_loader.current_address[11] ),
    .A2(_2767_),
    .ZN(_2768_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5641_ (.A1(\soc.rom_loader.current_address[11] ),
    .A2(_2767_),
    .Z(_2769_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _5642_ (.A1(_2745_),
    .A2(_2768_),
    .A3(_2769_),
    .ZN(_0468_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5643_ (.A1(\soc.rom_loader.current_address[12] ),
    .A2(_2769_),
    .ZN(_2770_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5644_ (.A1(\soc.rom_loader.current_address[12] ),
    .A2(_2769_),
    .Z(_2771_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _5645_ (.A1(_2745_),
    .A2(_2770_),
    .A3(_2771_),
    .ZN(_0469_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5646_ (.A1(_2089_),
    .A2(\soc.rom_loader.was_loading ),
    .B1(_2771_),
    .B2(\soc.rom_loader.current_address[13] ),
    .ZN(_2772_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5647_ (.A1(\soc.rom_loader.current_address[13] ),
    .A2(_2771_),
    .B(_2772_),
    .ZN(_0470_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5648_ (.A1(\soc.rom_loader.current_address[13] ),
    .A2(_2771_),
    .ZN(_2773_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5649_ (.A1(\soc.rom_loader.current_address[14] ),
    .A2(_2773_),
    .Z(_2774_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5650_ (.A1(_2746_),
    .A2(_2774_),
    .ZN(_0471_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5651_ (.I(net45),
    .ZN(_2775_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5652_ (.A1(\soc.rom_loader.wait_fall_clk ),
    .A2(\soc.rom_loader.rom_request ),
    .B(_0175_),
    .ZN(_2776_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5653_ (.A1(\soc.rom_loader.wait_fall_clk ),
    .A2(_2775_),
    .B(_2776_),
    .ZN(_0472_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5654_ (.A1(_0846_),
    .A2(\soc.cpu.instruction[4] ),
    .ZN(_2777_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5655_ (.I(_2777_),
    .Z(_2778_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5656_ (.I(_2777_),
    .Z(_2779_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5657_ (.A1(\soc.cpu.ALU.x[0] ),
    .A2(_2779_),
    .ZN(_2780_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5658_ (.A1(_0878_),
    .A2(_2778_),
    .B(_2780_),
    .ZN(_0474_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5659_ (.A1(\soc.cpu.ALU.x[1] ),
    .A2(_2779_),
    .ZN(_2781_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5660_ (.A1(_0902_),
    .A2(_2778_),
    .B(_2781_),
    .ZN(_0475_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5661_ (.A1(\soc.cpu.ALU.x[2] ),
    .A2(_2779_),
    .ZN(_2782_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5662_ (.A1(_0920_),
    .A2(_2778_),
    .B(_2782_),
    .ZN(_0476_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5663_ (.A1(\soc.cpu.ALU.x[3] ),
    .A2(_2779_),
    .ZN(_2783_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5664_ (.A1(_0942_),
    .A2(_2778_),
    .B(_2783_),
    .ZN(_0477_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5665_ (.I(_2777_),
    .Z(_2784_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5666_ (.A1(\soc.cpu.ALU.x[4] ),
    .A2(_2784_),
    .ZN(_2785_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5667_ (.A1(_0958_),
    .A2(_2778_),
    .B(_2785_),
    .ZN(_0478_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5668_ (.A1(\soc.cpu.ALU.x[5] ),
    .A2(_2784_),
    .ZN(_2786_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5669_ (.A1(_0970_),
    .A2(_2778_),
    .B(_2786_),
    .ZN(_0479_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5670_ (.A1(\soc.cpu.ALU.x[6] ),
    .A2(_2784_),
    .ZN(_2787_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5671_ (.A1(_0989_),
    .A2(_2778_),
    .B(_2787_),
    .ZN(_0480_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5672_ (.A1(\soc.cpu.ALU.x[7] ),
    .A2(_2784_),
    .ZN(_2788_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5673_ (.A1(_1002_),
    .A2(_2778_),
    .B(_2788_),
    .ZN(_0481_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5674_ (.A1(\soc.cpu.ALU.x[8] ),
    .A2(_2784_),
    .ZN(_2789_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5675_ (.A1(_1024_),
    .A2(_2778_),
    .B(_2789_),
    .ZN(_0482_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5676_ (.A1(\soc.cpu.ALU.x[9] ),
    .A2(_2784_),
    .ZN(_2790_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5677_ (.A1(_1039_),
    .A2(_2778_),
    .B(_2790_),
    .ZN(_0483_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5678_ (.A1(\soc.cpu.ALU.x[10] ),
    .A2(_2784_),
    .ZN(_2791_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5679_ (.A1(_1058_),
    .A2(_2779_),
    .B(_2791_),
    .ZN(_0484_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5680_ (.A1(\soc.cpu.ALU.x[11] ),
    .A2(_2784_),
    .ZN(_2792_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5681_ (.A1(_1069_),
    .A2(_2779_),
    .B(_2792_),
    .ZN(_0485_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5682_ (.A1(\soc.cpu.ALU.x[12] ),
    .A2(_2784_),
    .ZN(_2793_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5683_ (.A1(_1092_),
    .A2(_2779_),
    .B(_2793_),
    .ZN(_0486_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5684_ (.A1(\soc.cpu.ALU.x[13] ),
    .A2(_2784_),
    .ZN(_2794_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5685_ (.A1(_1108_),
    .A2(_2779_),
    .B(_2794_),
    .ZN(_0487_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5686_ (.A1(\soc.cpu.ALU.x[14] ),
    .A2(_2777_),
    .ZN(_2795_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5687_ (.A1(_1123_),
    .A2(_2779_),
    .B(_2795_),
    .ZN(_0488_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5688_ (.A1(\soc.cpu.ALU.x[15] ),
    .A2(_2777_),
    .ZN(_2796_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5689_ (.A1(_1669_),
    .A2(_2779_),
    .B(_2796_),
    .ZN(_0489_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _5690_ (.A1(_0700_),
    .A2(_2703_),
    .A3(_0698_),
    .ZN(_2797_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _5691_ (.I(_2797_),
    .Z(_2798_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _5692_ (.I(_2798_),
    .Z(_2799_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5693_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[6][0] ),
    .I1(\soc.spi_video_ram_1.fifo_in_data[0] ),
    .S(_2799_),
    .Z(_2800_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5694_ (.I(_2800_),
    .Z(_0490_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5695_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[6][1] ),
    .I1(\soc.spi_video_ram_1.fifo_in_data[1] ),
    .S(_2799_),
    .Z(_2801_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5696_ (.I(_2801_),
    .Z(_0491_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5697_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[6][2] ),
    .I1(\soc.spi_video_ram_1.fifo_in_data[2] ),
    .S(_2799_),
    .Z(_2802_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5698_ (.I(_2802_),
    .Z(_0492_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5699_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[6][3] ),
    .I1(\soc.spi_video_ram_1.fifo_in_data[3] ),
    .S(_2799_),
    .Z(_2803_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5700_ (.I(_2803_),
    .Z(_0493_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5701_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[6][4] ),
    .I1(\soc.spi_video_ram_1.fifo_in_data[4] ),
    .S(_2799_),
    .Z(_2804_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5702_ (.I(_2804_),
    .Z(_0494_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5703_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[6][5] ),
    .I1(\soc.spi_video_ram_1.fifo_in_data[5] ),
    .S(_2799_),
    .Z(_2805_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5704_ (.I(_2805_),
    .Z(_0495_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5705_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[6][6] ),
    .I1(\soc.spi_video_ram_1.fifo_in_data[6] ),
    .S(_2799_),
    .Z(_2806_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5706_ (.I(_2806_),
    .Z(_0496_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5707_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[6][7] ),
    .I1(\soc.spi_video_ram_1.fifo_in_data[7] ),
    .S(_2799_),
    .Z(_2807_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5708_ (.I(_2807_),
    .Z(_0497_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5709_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[6][8] ),
    .I1(\soc.spi_video_ram_1.fifo_in_data[8] ),
    .S(_2799_),
    .Z(_2808_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5710_ (.I(_2808_),
    .Z(_0498_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5711_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[6][9] ),
    .I1(\soc.spi_video_ram_1.fifo_in_data[9] ),
    .S(_2799_),
    .Z(_2809_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5712_ (.I(_2809_),
    .Z(_0499_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _5713_ (.I(_2797_),
    .Z(_2810_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5714_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[6][10] ),
    .I1(\soc.spi_video_ram_1.fifo_in_data[10] ),
    .S(_2810_),
    .Z(_2811_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5715_ (.I(_2811_),
    .Z(_0500_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5716_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[6][11] ),
    .I1(\soc.spi_video_ram_1.fifo_in_data[11] ),
    .S(_2810_),
    .Z(_2812_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5717_ (.I(_2812_),
    .Z(_0501_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5718_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[6][12] ),
    .I1(\soc.spi_video_ram_1.fifo_in_data[12] ),
    .S(_2810_),
    .Z(_2813_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5719_ (.I(_2813_),
    .Z(_0502_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5720_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[6][13] ),
    .I1(\soc.spi_video_ram_1.fifo_in_data[13] ),
    .S(_2810_),
    .Z(_2814_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5721_ (.I(_2814_),
    .Z(_0503_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5722_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[6][14] ),
    .I1(\soc.spi_video_ram_1.fifo_in_data[14] ),
    .S(_2810_),
    .Z(_2815_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5723_ (.I(_2815_),
    .Z(_0504_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5724_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[6][15] ),
    .I1(\soc.spi_video_ram_1.fifo_in_data[15] ),
    .S(_2810_),
    .Z(_2816_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5725_ (.I(_2816_),
    .Z(_0505_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5726_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[6][16] ),
    .I1(\soc.spi_video_ram_1.fifo_in_address[0] ),
    .S(_2810_),
    .Z(_2817_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5727_ (.I(_2817_),
    .Z(_0506_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5728_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[6][17] ),
    .I1(\soc.spi_video_ram_1.fifo_in_address[1] ),
    .S(_2810_),
    .Z(_2818_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5729_ (.I(_2818_),
    .Z(_0507_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5730_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[6][18] ),
    .I1(\soc.spi_video_ram_1.fifo_in_address[2] ),
    .S(_2810_),
    .Z(_2819_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5731_ (.I(_2819_),
    .Z(_0508_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5732_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[6][19] ),
    .I1(\soc.spi_video_ram_1.fifo_in_address[3] ),
    .S(_2810_),
    .Z(_2820_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5733_ (.I(_2820_),
    .Z(_0509_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5734_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[6][20] ),
    .I1(\soc.spi_video_ram_1.fifo_in_address[4] ),
    .S(_2798_),
    .Z(_2821_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5735_ (.I(_2821_),
    .Z(_0510_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5736_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[6][21] ),
    .I1(\soc.spi_video_ram_1.fifo_in_address[5] ),
    .S(_2798_),
    .Z(_2822_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5737_ (.I(_2822_),
    .Z(_0511_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5738_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[6][22] ),
    .I1(\soc.spi_video_ram_1.fifo_in_address[6] ),
    .S(_2798_),
    .Z(_2823_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5739_ (.I(_2823_),
    .Z(_0512_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5740_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[6][23] ),
    .I1(\soc.spi_video_ram_1.fifo_in_address[7] ),
    .S(_2798_),
    .Z(_2824_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5741_ (.I(_2824_),
    .Z(_0513_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5742_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[6][24] ),
    .I1(\soc.spi_video_ram_1.fifo_in_address[8] ),
    .S(_2798_),
    .Z(_2825_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5743_ (.I(_2825_),
    .Z(_0514_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5744_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[6][25] ),
    .I1(\soc.spi_video_ram_1.fifo_in_address[9] ),
    .S(_2798_),
    .Z(_2826_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5745_ (.I(_2826_),
    .Z(_0515_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5746_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[6][26] ),
    .I1(\soc.spi_video_ram_1.fifo_in_address[10] ),
    .S(_2798_),
    .Z(_2827_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5747_ (.I(_2827_),
    .Z(_0516_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5748_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[6][27] ),
    .I1(\soc.spi_video_ram_1.fifo_in_address[11] ),
    .S(_2798_),
    .Z(_2828_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5749_ (.I(_2828_),
    .Z(_0517_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5750_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[6][28] ),
    .I1(\soc.spi_video_ram_1.fifo_in_address[12] ),
    .S(_2798_),
    .Z(_2829_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5751_ (.I(_2829_),
    .Z(_0518_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5752_ (.A1(_0689_),
    .A2(_2690_),
    .ZN(_2830_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5753_ (.I(_2830_),
    .Z(_0535_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5754_ (.A1(net84),
    .A2(_0535_),
    .ZN(_2831_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5755_ (.A1(net84),
    .A2(_2691_),
    .B(_2831_),
    .ZN(_0519_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5756_ (.A1(_0922_),
    .A2(_1038_),
    .Z(_2832_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5757_ (.A1(_0922_),
    .A2(_1057_),
    .Z(_2833_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5758_ (.A1(_0990_),
    .A2(_1091_),
    .Z(_2834_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _5759_ (.A1(_0878_),
    .A2(_0902_),
    .A3(_0920_),
    .A4(_0942_),
    .Z(_2835_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _5760_ (.A1(_0958_),
    .A2(_0970_),
    .A3(_1002_),
    .A4(_2835_),
    .Z(_2836_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5761_ (.A1(_0989_),
    .A2(_1024_),
    .A3(_2836_),
    .ZN(_2837_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _5762_ (.A1(_2832_),
    .A2(_2833_),
    .A3(_2834_),
    .A4(_2837_),
    .ZN(_2838_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _5763_ (.A1(_1069_),
    .A2(_1108_),
    .A3(_2838_),
    .Z(_2839_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5764_ (.A1(_1123_),
    .A2(_2839_),
    .B(_0847_),
    .ZN(_2840_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5765_ (.I(\soc.cpu.DMuxJMP.sel[1] ),
    .ZN(_2841_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5766_ (.A1(_0990_),
    .A2(_1122_),
    .Z(_2842_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5767_ (.A1(_1069_),
    .A2(_1108_),
    .A3(_2838_),
    .ZN(_2843_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _5768_ (.A1(_2841_),
    .A2(_2842_),
    .A3(_2843_),
    .B(_1669_),
    .ZN(_2844_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _5769_ (.A1(\soc.cpu.DMuxJMP.sel[2] ),
    .A2(_1669_),
    .B1(_2840_),
    .B2(_2844_),
    .C(_0846_),
    .ZN(_2845_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5770_ (.I(_2845_),
    .Z(_2846_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5771_ (.I(_2845_),
    .Z(_2847_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5772_ (.A1(\soc.cpu.PC.in[0] ),
    .A2(_2847_),
    .ZN(_2848_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5773_ (.I(_0743_),
    .Z(_2849_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _5774_ (.A1(\soc.cpu.PC.REG.data[0] ),
    .A2(_2846_),
    .B(_2848_),
    .C(_2849_),
    .ZN(_0520_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5775_ (.A1(\soc.cpu.PC.REG.data[0] ),
    .A2(\soc.cpu.PC.REG.data[1] ),
    .ZN(_2850_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5776_ (.I(_2845_),
    .Z(_2851_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5777_ (.A1(\soc.cpu.PC.in[1] ),
    .A2(_2851_),
    .ZN(_2852_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _5778_ (.A1(_2846_),
    .A2(_2850_),
    .B(_2852_),
    .C(_2849_),
    .ZN(_0521_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5779_ (.A1(\soc.cpu.PC.REG.data[0] ),
    .A2(\soc.cpu.PC.REG.data[1] ),
    .ZN(_2853_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5780_ (.A1(\soc.cpu.PC.REG.data[2] ),
    .A2(_2853_),
    .Z(_2854_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5781_ (.A1(\soc.cpu.PC.in[2] ),
    .A2(_2851_),
    .ZN(_2855_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _5782_ (.A1(_2846_),
    .A2(_2854_),
    .B(_2855_),
    .C(_2849_),
    .ZN(_0522_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5783_ (.A1(\soc.cpu.PC.REG.data[0] ),
    .A2(\soc.cpu.PC.REG.data[1] ),
    .A3(\soc.cpu.PC.REG.data[2] ),
    .ZN(_2856_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5784_ (.A1(\soc.cpu.PC.REG.data[3] ),
    .A2(_2856_),
    .Z(_2857_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5785_ (.A1(\soc.cpu.PC.in[3] ),
    .A2(_2851_),
    .ZN(_2858_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _5786_ (.A1(_2846_),
    .A2(_2857_),
    .B(_2858_),
    .C(_2849_),
    .ZN(_0523_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5787_ (.A1(_2300_),
    .A2(_2856_),
    .ZN(_2859_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5788_ (.A1(\soc.cpu.PC.REG.data[4] ),
    .A2(_2859_),
    .ZN(_2860_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5789_ (.I(_2531_),
    .Z(_2861_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5790_ (.A1(\soc.cpu.PC.in[4] ),
    .A2(_2847_),
    .B(_2861_),
    .ZN(_2862_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5791_ (.A1(_2846_),
    .A2(_2860_),
    .B(_2862_),
    .ZN(_0524_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5792_ (.A1(\soc.cpu.PC.REG.data[4] ),
    .A2(_2859_),
    .Z(_2863_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5793_ (.A1(\soc.cpu.PC.REG.data[5] ),
    .A2(_2863_),
    .ZN(_2864_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5794_ (.A1(\soc.cpu.PC.in[5] ),
    .A2(_2847_),
    .B(_2861_),
    .ZN(_2865_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5795_ (.A1(_2846_),
    .A2(_2864_),
    .B(_2865_),
    .ZN(_0525_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5796_ (.A1(\soc.cpu.PC.REG.data[5] ),
    .A2(_2863_),
    .ZN(_2866_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5797_ (.A1(\soc.cpu.PC.REG.data[6] ),
    .A2(_2866_),
    .Z(_2867_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5798_ (.A1(\soc.cpu.PC.in[6] ),
    .A2(_2847_),
    .B(_2861_),
    .ZN(_2868_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5799_ (.A1(_2846_),
    .A2(_2867_),
    .B(_2868_),
    .ZN(_0526_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5800_ (.A1(\soc.cpu.PC.REG.data[5] ),
    .A2(\soc.cpu.PC.REG.data[6] ),
    .A3(_2863_),
    .ZN(_2869_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5801_ (.A1(\soc.cpu.PC.REG.data[7] ),
    .A2(_2869_),
    .Z(_2870_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5802_ (.A1(\soc.cpu.PC.in[7] ),
    .A2(_2851_),
    .ZN(_2871_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _5803_ (.A1(_2846_),
    .A2(_2870_),
    .B(_2871_),
    .C(_2849_),
    .ZN(_0527_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5804_ (.A1(_2310_),
    .A2(_2869_),
    .ZN(_2872_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5805_ (.A1(\soc.cpu.PC.REG.data[8] ),
    .A2(_2872_),
    .ZN(_2873_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5806_ (.A1(\soc.cpu.PC.in[8] ),
    .A2(_2851_),
    .ZN(_2874_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _5807_ (.A1(_2846_),
    .A2(_2873_),
    .B(_2874_),
    .C(_2849_),
    .ZN(_0528_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5808_ (.A1(\soc.cpu.PC.REG.data[8] ),
    .A2(_2872_),
    .ZN(_2875_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5809_ (.A1(\soc.cpu.PC.REG.data[9] ),
    .A2(_2875_),
    .Z(_2876_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5810_ (.A1(\soc.cpu.PC.in[9] ),
    .A2(_2851_),
    .ZN(_2877_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _5811_ (.A1(_2847_),
    .A2(_2876_),
    .B(_2877_),
    .C(_2849_),
    .ZN(_0529_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5812_ (.A1(\soc.cpu.PC.REG.data[8] ),
    .A2(\soc.cpu.PC.REG.data[9] ),
    .A3(_2872_),
    .ZN(_2878_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5813_ (.A1(\soc.cpu.PC.REG.data[10] ),
    .A2(_2878_),
    .Z(_2879_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5814_ (.A1(\soc.cpu.PC.in[10] ),
    .A2(_2851_),
    .ZN(_2880_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _5815_ (.A1(_2847_),
    .A2(_2879_),
    .B(_2880_),
    .C(_2849_),
    .ZN(_0530_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5816_ (.A1(_2318_),
    .A2(_2878_),
    .ZN(_2881_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5817_ (.A1(\soc.cpu.PC.REG.data[11] ),
    .A2(_2881_),
    .ZN(_2882_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5818_ (.A1(\soc.cpu.PC.in[11] ),
    .A2(_2847_),
    .B(_2861_),
    .ZN(_2883_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5819_ (.A1(_2846_),
    .A2(_2882_),
    .B(_2883_),
    .ZN(_0531_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5820_ (.A1(\soc.cpu.PC.REG.data[11] ),
    .A2(_2881_),
    .ZN(_2884_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5821_ (.A1(\soc.cpu.PC.REG.data[12] ),
    .A2(_2884_),
    .Z(_2885_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5822_ (.A1(\soc.cpu.PC.in[12] ),
    .A2(_2851_),
    .ZN(_2886_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _5823_ (.A1(_2847_),
    .A2(_2885_),
    .B(_2886_),
    .C(_2849_),
    .ZN(_0532_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5824_ (.A1(\soc.cpu.PC.REG.data[11] ),
    .A2(\soc.cpu.PC.REG.data[12] ),
    .A3(_2881_),
    .ZN(_2887_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5825_ (.A1(\soc.cpu.PC.REG.data[13] ),
    .A2(_2887_),
    .Z(_2888_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5826_ (.A1(\soc.cpu.PC.in[13] ),
    .A2(_2851_),
    .ZN(_2889_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _5827_ (.A1(_2847_),
    .A2(_2888_),
    .B(_2889_),
    .C(_2849_),
    .ZN(_0533_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _5828_ (.A1(\soc.cpu.PC.REG.data[11] ),
    .A2(\soc.cpu.PC.REG.data[12] ),
    .A3(\soc.cpu.PC.REG.data[13] ),
    .A4(_2881_),
    .ZN(_2890_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5829_ (.A1(\soc.cpu.PC.REG.data[14] ),
    .A2(_2890_),
    .Z(_2891_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5830_ (.A1(\soc.cpu.PC.in[14] ),
    .A2(_2851_),
    .ZN(_2892_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _5831_ (.A1(_2847_),
    .A2(_2891_),
    .B(_2892_),
    .C(_0743_),
    .ZN(_0534_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5832_ (.A1(_2688_),
    .A2(_2689_),
    .A3(_2692_),
    .ZN(_2893_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5833_ (.A1(net85),
    .A2(_2893_),
    .Z(_2894_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5834_ (.A1(_0744_),
    .A2(_2894_),
    .Z(_2895_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5835_ (.I(_2895_),
    .Z(_2896_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5836_ (.I(_2896_),
    .Z(_2897_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5837_ (.I(net85),
    .ZN(_2898_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5838_ (.A1(_2898_),
    .A2(\soc.hack_clk_strobe ),
    .A3(_2893_),
    .ZN(_2899_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5839_ (.A1(\soc.synch_hack_writeM ),
    .A2(_2899_),
    .ZN(_2900_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5840_ (.A1(_2897_),
    .A2(_2900_),
    .ZN(_0536_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5841_ (.A1(_2896_),
    .A2(_2899_),
    .ZN(_2901_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _5842_ (.I(_2901_),
    .Z(_2902_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _5843_ (.I(_2902_),
    .Z(_2903_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5844_ (.A1(\soc.ram_encoder_0.address[0] ),
    .A2(_2903_),
    .ZN(_2904_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5845_ (.A1(_0855_),
    .A2(_2903_),
    .B(_2904_),
    .ZN(_0537_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5846_ (.I0(\soc.ram_encoder_0.address[1] ),
    .I1(\soc.cpu.AReg.data[1] ),
    .S(_2903_),
    .Z(_2905_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5847_ (.I(_2905_),
    .Z(_0538_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5848_ (.A1(\soc.ram_encoder_0.address[2] ),
    .A2(_2903_),
    .ZN(_2906_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5849_ (.A1(_0908_),
    .A2(_2903_),
    .B(_2906_),
    .ZN(_0539_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5850_ (.I0(\soc.ram_encoder_0.address[3] ),
    .I1(\soc.cpu.AReg.data[3] ),
    .S(_2903_),
    .Z(_2907_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5851_ (.I(_2907_),
    .Z(_0540_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5852_ (.I0(\soc.ram_encoder_0.address[4] ),
    .I1(\soc.cpu.AReg.data[4] ),
    .S(_2903_),
    .Z(_2908_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5853_ (.I(_2908_),
    .Z(_0541_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5854_ (.I0(\soc.ram_encoder_0.address[5] ),
    .I1(\soc.cpu.AReg.data[5] ),
    .S(_2903_),
    .Z(_2909_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5855_ (.I(_2909_),
    .Z(_0542_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5856_ (.I0(\soc.ram_encoder_0.address[6] ),
    .I1(\soc.cpu.AReg.data[6] ),
    .S(_2902_),
    .Z(_2910_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5857_ (.I(_2910_),
    .Z(_0543_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5858_ (.I0(\soc.ram_encoder_0.address[7] ),
    .I1(\soc.cpu.AReg.data[7] ),
    .S(_2902_),
    .Z(_2911_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5859_ (.I(_2911_),
    .Z(_0544_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5860_ (.I0(\soc.ram_encoder_0.address[8] ),
    .I1(\soc.cpu.AReg.data[8] ),
    .S(_2902_),
    .Z(_2912_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5861_ (.I(_2912_),
    .Z(_0545_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5862_ (.I0(\soc.ram_encoder_0.address[9] ),
    .I1(\soc.cpu.AReg.data[9] ),
    .S(_2902_),
    .Z(_2913_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5863_ (.I(_2913_),
    .Z(_0546_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5864_ (.I0(\soc.ram_encoder_0.address[10] ),
    .I1(\soc.cpu.AReg.data[10] ),
    .S(_2902_),
    .Z(_2914_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5865_ (.I(_2914_),
    .Z(_0547_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5866_ (.I0(\soc.ram_encoder_0.address[11] ),
    .I1(\soc.cpu.AReg.data[11] ),
    .S(_2902_),
    .Z(_2915_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5867_ (.I(_2915_),
    .Z(_0548_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5868_ (.I0(\soc.ram_encoder_0.address[12] ),
    .I1(\soc.cpu.AReg.data[12] ),
    .S(_2902_),
    .Z(_2916_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5869_ (.I(_2916_),
    .Z(_0549_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5870_ (.A1(\soc.ram_encoder_0.address[13] ),
    .A2(_2903_),
    .ZN(_2917_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5871_ (.A1(_0745_),
    .A2(_2903_),
    .B(_2917_),
    .ZN(_0550_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5872_ (.I0(\soc.ram_encoder_0.address[14] ),
    .I1(\soc.cpu.AReg.data[14] ),
    .S(_2902_),
    .Z(_2918_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5873_ (.I(_2918_),
    .Z(_0551_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5874_ (.I(_2899_),
    .ZN(_0552_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5875_ (.I(_2897_),
    .ZN(_0553_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5876_ (.A1(_2898_),
    .A2(\soc.hack_clk_strobe ),
    .ZN(_2919_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5877_ (.A1(_2738_),
    .A2(_2919_),
    .ZN(_0554_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5878_ (.A1(_2293_),
    .A2(net45),
    .B(\soc.boot_loading_offset[0] ),
    .ZN(_2920_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5879_ (.A1(_1209_),
    .A2(_2739_),
    .ZN(_2921_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _5880_ (.A1(_1461_),
    .A2(_2920_),
    .A3(_2921_),
    .ZN(_0555_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5881_ (.A1(\soc.boot_loading_offset[1] ),
    .A2(_2921_),
    .B(_0689_),
    .ZN(_2922_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5882_ (.A1(\soc.boot_loading_offset[1] ),
    .A2(_2921_),
    .B(_2922_),
    .ZN(_2923_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5883_ (.I(_2923_),
    .ZN(_0556_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5884_ (.A1(\soc.boot_loading_offset[1] ),
    .A2(_2921_),
    .B(\soc.boot_loading_offset[2] ),
    .ZN(_2924_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _5885_ (.A1(\soc.boot_loading_offset[2] ),
    .A2(\soc.boot_loading_offset[1] ),
    .A3(_2921_),
    .Z(_2925_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _5886_ (.A1(_1461_),
    .A2(_2924_),
    .A3(_2925_),
    .ZN(_0557_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5887_ (.A1(\soc.boot_loading_offset[3] ),
    .A2(_2925_),
    .B(_0675_),
    .ZN(_2926_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5888_ (.A1(\soc.boot_loading_offset[3] ),
    .A2(_2925_),
    .B(_2926_),
    .ZN(_0558_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5889_ (.A1(\soc.boot_loading_offset[3] ),
    .A2(_2925_),
    .ZN(_2927_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5890_ (.A1(\soc.boot_loading_offset[4] ),
    .A2(_2927_),
    .Z(_2928_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5891_ (.A1(_2471_),
    .A2(_2928_),
    .ZN(_0559_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5892_ (.A1(net85),
    .A2(\soc.hack_clk_strobe ),
    .ZN(_2929_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5893_ (.I(net19),
    .ZN(_2930_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5894_ (.A1(_2861_),
    .A2(_2929_),
    .B(_2930_),
    .ZN(_0560_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5895_ (.A1(\soc.hack_wait_clocks[0] ),
    .A2(_2929_),
    .ZN(_2931_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5896_ (.A1(\soc.hack_wait_clocks[0] ),
    .A2(_2929_),
    .ZN(_2932_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5897_ (.A1(\soc.hack_wait_clocks[1] ),
    .A2(_2932_),
    .ZN(_2933_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5898_ (.A1(_2931_),
    .A2(_2933_),
    .B(_0741_),
    .ZN(_0561_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5899_ (.I(\soc.hack_wait_clocks[1] ),
    .ZN(_2934_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5900_ (.I(_0741_),
    .ZN(_2935_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5901_ (.A1(_2934_),
    .A2(_2932_),
    .B(_2935_),
    .ZN(_0562_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _5902_ (.A1(\soc.cpu.AReg.data[0] ),
    .A2(_0744_),
    .A3(_0864_),
    .A4(_0930_),
    .ZN(_2936_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5903_ (.A1(net77),
    .A2(_2936_),
    .B(_2861_),
    .ZN(_2937_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5904_ (.A1(_0878_),
    .A2(_2936_),
    .B(_2937_),
    .ZN(_0563_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5905_ (.A1(net78),
    .A2(_2936_),
    .B(_2861_),
    .ZN(_2938_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5906_ (.A1(_0902_),
    .A2(_2936_),
    .B(_2938_),
    .ZN(_0564_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5907_ (.A1(net79),
    .A2(_2936_),
    .B(_2861_),
    .ZN(_2939_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5908_ (.A1(_0920_),
    .A2(_2936_),
    .B(_2939_),
    .ZN(_0565_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5909_ (.A1(net80),
    .A2(_2936_),
    .B(_2861_),
    .ZN(_2940_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5910_ (.A1(_0942_),
    .A2(_2936_),
    .B(_2940_),
    .ZN(_0566_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5911_ (.I(net14),
    .ZN(_2941_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5912_ (.A1(_0744_),
    .A2(_0867_),
    .Z(_2942_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5913_ (.I(_2942_),
    .Z(_2943_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5914_ (.A1(\soc.gpio_i_stored[0] ),
    .A2(_2943_),
    .B(_2861_),
    .ZN(_2944_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5915_ (.A1(_2941_),
    .A2(_2943_),
    .B(_2944_),
    .ZN(_0567_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5916_ (.I(net15),
    .ZN(_2945_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5917_ (.A1(\soc.gpio_i_stored[1] ),
    .A2(_2943_),
    .B(_2531_),
    .ZN(_2946_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5918_ (.A1(_2945_),
    .A2(_2943_),
    .B(_2946_),
    .ZN(_0568_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5919_ (.I(net16),
    .ZN(_2947_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5920_ (.A1(\soc.gpio_i_stored[2] ),
    .A2(_2943_),
    .B(_2531_),
    .ZN(_2948_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5921_ (.A1(_2947_),
    .A2(_2943_),
    .B(_2948_),
    .ZN(_0569_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5922_ (.I(net17),
    .ZN(_2949_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5923_ (.A1(\soc.gpio_i_stored[3] ),
    .A2(_2943_),
    .B(_2531_),
    .ZN(_2950_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5924_ (.A1(_2949_),
    .A2(_2943_),
    .B(_2950_),
    .ZN(_0570_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _5925_ (.A1(\soc.spi_video_ram_1.write_fifo.write_pointer[2] ),
    .A2(_0694_),
    .A3(_0698_),
    .ZN(_2951_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _5926_ (.I(_2951_),
    .Z(_2952_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _5927_ (.I(_2952_),
    .Z(_2953_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5928_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[0][0] ),
    .I1(\soc.spi_video_ram_1.fifo_in_data[0] ),
    .S(_2953_),
    .Z(_2954_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5929_ (.I(_2954_),
    .Z(_0571_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5930_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[0][1] ),
    .I1(\soc.spi_video_ram_1.fifo_in_data[1] ),
    .S(_2953_),
    .Z(_2955_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5931_ (.I(_2955_),
    .Z(_0572_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5932_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[0][2] ),
    .I1(\soc.spi_video_ram_1.fifo_in_data[2] ),
    .S(_2953_),
    .Z(_2956_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5933_ (.I(_2956_),
    .Z(_0573_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5934_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[0][3] ),
    .I1(\soc.spi_video_ram_1.fifo_in_data[3] ),
    .S(_2953_),
    .Z(_2957_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5935_ (.I(_2957_),
    .Z(_0574_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5936_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[0][4] ),
    .I1(\soc.spi_video_ram_1.fifo_in_data[4] ),
    .S(_2953_),
    .Z(_2958_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5937_ (.I(_2958_),
    .Z(_0575_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5938_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[0][5] ),
    .I1(\soc.spi_video_ram_1.fifo_in_data[5] ),
    .S(_2953_),
    .Z(_2959_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5939_ (.I(_2959_),
    .Z(_0576_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5940_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[0][6] ),
    .I1(\soc.spi_video_ram_1.fifo_in_data[6] ),
    .S(_2953_),
    .Z(_2960_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5941_ (.I(_2960_),
    .Z(_0577_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5942_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[0][7] ),
    .I1(\soc.spi_video_ram_1.fifo_in_data[7] ),
    .S(_2953_),
    .Z(_2961_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5943_ (.I(_2961_),
    .Z(_0578_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5944_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[0][8] ),
    .I1(\soc.spi_video_ram_1.fifo_in_data[8] ),
    .S(_2953_),
    .Z(_2962_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5945_ (.I(_2962_),
    .Z(_0579_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5946_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[0][9] ),
    .I1(\soc.spi_video_ram_1.fifo_in_data[9] ),
    .S(_2953_),
    .Z(_2963_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5947_ (.I(_2963_),
    .Z(_0580_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _5948_ (.I(_2951_),
    .Z(_2964_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5949_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[0][10] ),
    .I1(\soc.spi_video_ram_1.fifo_in_data[10] ),
    .S(_2964_),
    .Z(_2965_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5950_ (.I(_2965_),
    .Z(_0581_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5951_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[0][11] ),
    .I1(\soc.spi_video_ram_1.fifo_in_data[11] ),
    .S(_2964_),
    .Z(_2966_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5952_ (.I(_2966_),
    .Z(_0582_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5953_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[0][12] ),
    .I1(\soc.spi_video_ram_1.fifo_in_data[12] ),
    .S(_2964_),
    .Z(_2967_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5954_ (.I(_2967_),
    .Z(_0583_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5955_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[0][13] ),
    .I1(\soc.spi_video_ram_1.fifo_in_data[13] ),
    .S(_2964_),
    .Z(_2968_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5956_ (.I(_2968_),
    .Z(_0584_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5957_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[0][14] ),
    .I1(\soc.spi_video_ram_1.fifo_in_data[14] ),
    .S(_2964_),
    .Z(_2969_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5958_ (.I(_2969_),
    .Z(_0585_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5959_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[0][15] ),
    .I1(\soc.spi_video_ram_1.fifo_in_data[15] ),
    .S(_2964_),
    .Z(_2970_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5960_ (.I(_2970_),
    .Z(_0586_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5961_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[0][16] ),
    .I1(\soc.spi_video_ram_1.fifo_in_address[0] ),
    .S(_2964_),
    .Z(_2971_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5962_ (.I(_2971_),
    .Z(_0587_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5963_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[0][17] ),
    .I1(\soc.spi_video_ram_1.fifo_in_address[1] ),
    .S(_2964_),
    .Z(_2972_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5964_ (.I(_2972_),
    .Z(_0588_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5965_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[0][18] ),
    .I1(\soc.spi_video_ram_1.fifo_in_address[2] ),
    .S(_2964_),
    .Z(_2973_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5966_ (.I(_2973_),
    .Z(_0589_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5967_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[0][19] ),
    .I1(\soc.spi_video_ram_1.fifo_in_address[3] ),
    .S(_2964_),
    .Z(_2974_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5968_ (.I(_2974_),
    .Z(_0590_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5969_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[0][20] ),
    .I1(\soc.spi_video_ram_1.fifo_in_address[4] ),
    .S(_2952_),
    .Z(_2975_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5970_ (.I(_2975_),
    .Z(_0591_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5971_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[0][21] ),
    .I1(\soc.spi_video_ram_1.fifo_in_address[5] ),
    .S(_2952_),
    .Z(_2976_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5972_ (.I(_2976_),
    .Z(_0592_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5973_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[0][22] ),
    .I1(\soc.spi_video_ram_1.fifo_in_address[6] ),
    .S(_2952_),
    .Z(_2977_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5974_ (.I(_2977_),
    .Z(_0593_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5975_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[0][23] ),
    .I1(\soc.spi_video_ram_1.fifo_in_address[7] ),
    .S(_2952_),
    .Z(_2978_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5976_ (.I(_2978_),
    .Z(_0594_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5977_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[0][24] ),
    .I1(\soc.spi_video_ram_1.fifo_in_address[8] ),
    .S(_2952_),
    .Z(_2979_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5978_ (.I(_2979_),
    .Z(_0595_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5979_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[0][25] ),
    .I1(\soc.spi_video_ram_1.fifo_in_address[9] ),
    .S(_2952_),
    .Z(_2980_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5980_ (.I(_2980_),
    .Z(_0596_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5981_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[0][26] ),
    .I1(\soc.spi_video_ram_1.fifo_in_address[10] ),
    .S(_2952_),
    .Z(_2981_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5982_ (.I(_2981_),
    .Z(_0597_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5983_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[0][27] ),
    .I1(\soc.spi_video_ram_1.fifo_in_address[11] ),
    .S(_2952_),
    .Z(_2982_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5984_ (.I(_2982_),
    .Z(_0598_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5985_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[0][28] ),
    .I1(\soc.spi_video_ram_1.fifo_in_address[12] ),
    .S(_2952_),
    .Z(_2983_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5986_ (.I(_2983_),
    .Z(_0599_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5987_ (.A1(_0700_),
    .A2(_2703_),
    .A3(_0698_),
    .ZN(_2984_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 _5988_ (.I(_2984_),
    .Z(_2985_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 _5989_ (.I(_2985_),
    .Z(_2986_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5990_ (.I0(\soc.spi_video_ram_1.fifo_in_data[0] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[1][0] ),
    .S(_2986_),
    .Z(_2987_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5991_ (.I(_2987_),
    .Z(_0600_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5992_ (.I(_2985_),
    .Z(_2988_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5993_ (.A1(\soc.spi_video_ram_1.fifo_in_data[1] ),
    .A2(_2988_),
    .ZN(_2989_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5994_ (.A1(_1698_),
    .A2(_2988_),
    .B(_2989_),
    .ZN(_0601_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5995_ (.I0(\soc.spi_video_ram_1.fifo_in_data[2] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[1][2] ),
    .S(_2986_),
    .Z(_2990_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5996_ (.I(_2990_),
    .Z(_0602_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5997_ (.I0(\soc.spi_video_ram_1.fifo_in_data[3] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[1][3] ),
    .S(_2986_),
    .Z(_2991_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5998_ (.I(_2991_),
    .Z(_0603_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5999_ (.I0(\soc.spi_video_ram_1.fifo_in_data[4] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[1][4] ),
    .S(_2986_),
    .Z(_2992_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6000_ (.I(_2992_),
    .Z(_0604_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6001_ (.A1(\soc.spi_video_ram_1.fifo_in_data[5] ),
    .A2(_2988_),
    .ZN(_2993_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6002_ (.A1(_1734_),
    .A2(_2988_),
    .B(_2993_),
    .ZN(_0605_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6003_ (.I0(\soc.spi_video_ram_1.fifo_in_data[6] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[1][6] ),
    .S(_2986_),
    .Z(_2994_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6004_ (.I(_2994_),
    .Z(_0606_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6005_ (.A1(\soc.spi_video_ram_1.fifo_in_data[7] ),
    .A2(_2988_),
    .ZN(_2995_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6006_ (.A1(_1775_),
    .A2(_2988_),
    .B(_2995_),
    .ZN(_0607_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6007_ (.A1(\soc.spi_video_ram_1.fifo_in_data[8] ),
    .A2(_2986_),
    .ZN(_2996_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6008_ (.A1(_1781_),
    .A2(_2988_),
    .B(_2996_),
    .ZN(_0608_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6009_ (.A1(\soc.spi_video_ram_1.fifo_in_data[9] ),
    .A2(_2986_),
    .ZN(_2997_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6010_ (.A1(_1799_),
    .A2(_2988_),
    .B(_2997_),
    .ZN(_0609_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6011_ (.I0(\soc.spi_video_ram_1.fifo_in_data[10] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[1][10] ),
    .S(_2986_),
    .Z(_2998_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6012_ (.I(_2998_),
    .Z(_0610_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _6013_ (.I(_2985_),
    .Z(_2999_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6014_ (.I0(\soc.spi_video_ram_1.fifo_in_data[11] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[1][11] ),
    .S(_2999_),
    .Z(_3000_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6015_ (.I(_3000_),
    .Z(_0611_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6016_ (.I0(\soc.spi_video_ram_1.fifo_in_data[12] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[1][12] ),
    .S(_2999_),
    .Z(_3001_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6017_ (.I(_3001_),
    .Z(_0612_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6018_ (.A1(\soc.spi_video_ram_1.fifo_in_data[13] ),
    .A2(_2986_),
    .ZN(_3002_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6019_ (.A1(_1860_),
    .A2(_2988_),
    .B(_3002_),
    .ZN(_0613_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6020_ (.A1(\soc.spi_video_ram_1.fifo_in_data[14] ),
    .A2(_2986_),
    .ZN(_3003_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6021_ (.A1(_1883_),
    .A2(_2988_),
    .B(_3003_),
    .ZN(_0614_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6022_ (.I0(\soc.spi_video_ram_1.fifo_in_data[15] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[1][15] ),
    .S(_2999_),
    .Z(_3004_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6023_ (.I(_3004_),
    .Z(_0615_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6024_ (.I0(\soc.spi_video_ram_1.fifo_in_address[0] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[1][16] ),
    .S(_2999_),
    .Z(_3005_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6025_ (.I(_3005_),
    .Z(_0616_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6026_ (.I0(\soc.spi_video_ram_1.fifo_in_address[1] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[1][17] ),
    .S(_2999_),
    .Z(_3006_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6027_ (.I(_3006_),
    .Z(_0617_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6028_ (.I0(\soc.spi_video_ram_1.fifo_in_address[2] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[1][18] ),
    .S(_2999_),
    .Z(_3007_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6029_ (.I(_3007_),
    .Z(_0618_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6030_ (.I0(\soc.spi_video_ram_1.fifo_in_address[3] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[1][19] ),
    .S(_2999_),
    .Z(_3008_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6031_ (.I(_3008_),
    .Z(_0619_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6032_ (.I0(\soc.spi_video_ram_1.fifo_in_address[4] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[1][20] ),
    .S(_2999_),
    .Z(_3009_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6033_ (.I(_3009_),
    .Z(_0620_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6034_ (.I0(\soc.spi_video_ram_1.fifo_in_address[5] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[1][21] ),
    .S(_2999_),
    .Z(_3010_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6035_ (.I(_3010_),
    .Z(_0621_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6036_ (.I0(\soc.spi_video_ram_1.fifo_in_address[6] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[1][22] ),
    .S(_2999_),
    .Z(_3011_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6037_ (.I(_3011_),
    .Z(_0622_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6038_ (.I0(\soc.spi_video_ram_1.fifo_in_address[7] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[1][23] ),
    .S(_2985_),
    .Z(_3012_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6039_ (.I(_3012_),
    .Z(_0623_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6040_ (.I0(\soc.spi_video_ram_1.fifo_in_address[8] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[1][24] ),
    .S(_2985_),
    .Z(_3013_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6041_ (.I(_3013_),
    .Z(_0624_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6042_ (.I0(\soc.spi_video_ram_1.fifo_in_address[9] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[1][25] ),
    .S(_2985_),
    .Z(_3014_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6043_ (.I(_3014_),
    .Z(_0625_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6044_ (.I0(\soc.spi_video_ram_1.fifo_in_address[10] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[1][26] ),
    .S(_2985_),
    .Z(_3015_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6045_ (.I(_3015_),
    .Z(_0626_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6046_ (.I0(\soc.spi_video_ram_1.fifo_in_address[11] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[1][27] ),
    .S(_2985_),
    .Z(_3016_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6047_ (.I(_3016_),
    .Z(_0627_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6048_ (.I0(\soc.spi_video_ram_1.fifo_in_address[12] ),
    .I1(\soc.spi_video_ram_1.write_fifo.fifo_mem[1][28] ),
    .S(_2985_),
    .Z(_3017_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6049_ (.I(_3017_),
    .Z(_0628_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _6050_ (.A1(\soc.spi_video_ram_1.write_fifo.write_pointer[2] ),
    .A2(_2703_),
    .A3(_0698_),
    .ZN(_3018_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _6051_ (.I(_3018_),
    .Z(_3019_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _6052_ (.I(_3019_),
    .Z(_3020_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6053_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[2][0] ),
    .I1(\soc.spi_video_ram_1.fifo_in_data[0] ),
    .S(_3020_),
    .Z(_3021_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6054_ (.I(_3021_),
    .Z(_0629_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6055_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[2][1] ),
    .I1(\soc.spi_video_ram_1.fifo_in_data[1] ),
    .S(_3020_),
    .Z(_3022_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6056_ (.I(_3022_),
    .Z(_0630_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6057_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[2][2] ),
    .I1(\soc.spi_video_ram_1.fifo_in_data[2] ),
    .S(_3020_),
    .Z(_3023_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6058_ (.I(_3023_),
    .Z(_0631_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6059_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[2][3] ),
    .I1(\soc.spi_video_ram_1.fifo_in_data[3] ),
    .S(_3020_),
    .Z(_3024_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6060_ (.I(_3024_),
    .Z(_0632_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6061_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[2][4] ),
    .I1(\soc.spi_video_ram_1.fifo_in_data[4] ),
    .S(_3020_),
    .Z(_3025_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6062_ (.I(_3025_),
    .Z(_0633_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6063_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[2][5] ),
    .I1(\soc.spi_video_ram_1.fifo_in_data[5] ),
    .S(_3020_),
    .Z(_3026_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6064_ (.I(_3026_),
    .Z(_0634_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6065_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[2][6] ),
    .I1(\soc.spi_video_ram_1.fifo_in_data[6] ),
    .S(_3020_),
    .Z(_3027_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6066_ (.I(_3027_),
    .Z(_0635_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6067_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[2][7] ),
    .I1(\soc.spi_video_ram_1.fifo_in_data[7] ),
    .S(_3020_),
    .Z(_3028_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6068_ (.I(_3028_),
    .Z(_0636_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6069_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[2][8] ),
    .I1(\soc.spi_video_ram_1.fifo_in_data[8] ),
    .S(_3020_),
    .Z(_3029_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6070_ (.I(_3029_),
    .Z(_0637_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6071_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[2][9] ),
    .I1(\soc.spi_video_ram_1.fifo_in_data[9] ),
    .S(_3020_),
    .Z(_3030_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6072_ (.I(_3030_),
    .Z(_0638_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _6073_ (.I(_3018_),
    .Z(_3031_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6074_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[2][10] ),
    .I1(\soc.spi_video_ram_1.fifo_in_data[10] ),
    .S(_3031_),
    .Z(_3032_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6075_ (.I(_3032_),
    .Z(_0639_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6076_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[2][11] ),
    .I1(\soc.spi_video_ram_1.fifo_in_data[11] ),
    .S(_3031_),
    .Z(_3033_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6077_ (.I(_3033_),
    .Z(_0640_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6078_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[2][12] ),
    .I1(\soc.spi_video_ram_1.fifo_in_data[12] ),
    .S(_3031_),
    .Z(_3034_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6079_ (.I(_3034_),
    .Z(_0641_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6080_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[2][13] ),
    .I1(\soc.spi_video_ram_1.fifo_in_data[13] ),
    .S(_3031_),
    .Z(_3035_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6081_ (.I(_3035_),
    .Z(_0642_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6082_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[2][14] ),
    .I1(\soc.spi_video_ram_1.fifo_in_data[14] ),
    .S(_3031_),
    .Z(_3036_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6083_ (.I(_3036_),
    .Z(_0643_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6084_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[2][15] ),
    .I1(\soc.spi_video_ram_1.fifo_in_data[15] ),
    .S(_3031_),
    .Z(_3037_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6085_ (.I(_3037_),
    .Z(_0644_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6086_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[2][16] ),
    .I1(\soc.spi_video_ram_1.fifo_in_address[0] ),
    .S(_3031_),
    .Z(_3038_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6087_ (.I(_3038_),
    .Z(_0645_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6088_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[2][17] ),
    .I1(\soc.spi_video_ram_1.fifo_in_address[1] ),
    .S(_3031_),
    .Z(_3039_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6089_ (.I(_3039_),
    .Z(_0646_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6090_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[2][18] ),
    .I1(\soc.spi_video_ram_1.fifo_in_address[2] ),
    .S(_3031_),
    .Z(_3040_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6091_ (.I(_3040_),
    .Z(_0647_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6092_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[2][19] ),
    .I1(\soc.spi_video_ram_1.fifo_in_address[3] ),
    .S(_3031_),
    .Z(_3041_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6093_ (.I(_3041_),
    .Z(_0648_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6094_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[2][20] ),
    .I1(\soc.spi_video_ram_1.fifo_in_address[4] ),
    .S(_3019_),
    .Z(_3042_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6095_ (.I(_3042_),
    .Z(_0649_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6096_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[2][21] ),
    .I1(\soc.spi_video_ram_1.fifo_in_address[5] ),
    .S(_3019_),
    .Z(_3043_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6097_ (.I(_3043_),
    .Z(_0650_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6098_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[2][22] ),
    .I1(\soc.spi_video_ram_1.fifo_in_address[6] ),
    .S(_3019_),
    .Z(_3044_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6099_ (.I(_3044_),
    .Z(_0651_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6100_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[2][23] ),
    .I1(\soc.spi_video_ram_1.fifo_in_address[7] ),
    .S(_3019_),
    .Z(_3045_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6101_ (.I(_3045_),
    .Z(_0652_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6102_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[2][24] ),
    .I1(\soc.spi_video_ram_1.fifo_in_address[8] ),
    .S(_3019_),
    .Z(_3046_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6103_ (.I(_3046_),
    .Z(_0653_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6104_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[2][25] ),
    .I1(\soc.spi_video_ram_1.fifo_in_address[9] ),
    .S(_3019_),
    .Z(_3047_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6105_ (.I(_3047_),
    .Z(_0654_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6106_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[2][26] ),
    .I1(\soc.spi_video_ram_1.fifo_in_address[10] ),
    .S(_3019_),
    .Z(_3048_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6107_ (.I(_3048_),
    .Z(_0655_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6108_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[2][27] ),
    .I1(\soc.spi_video_ram_1.fifo_in_address[11] ),
    .S(_3019_),
    .Z(_3049_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6109_ (.I(_3049_),
    .Z(_0656_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6110_ (.I0(\soc.spi_video_ram_1.write_fifo.fifo_mem[2][28] ),
    .I1(\soc.spi_video_ram_1.fifo_in_address[12] ),
    .S(_3019_),
    .Z(_3050_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6111_ (.I(_3050_),
    .Z(_0657_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _6112_ (.A1(_2894_),
    .A2(_2919_),
    .ZN(_3051_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _6113_ (.I(_3051_),
    .Z(_3052_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _6114_ (.A1(_0878_),
    .A2(_2897_),
    .B1(_3052_),
    .B2(_2541_),
    .ZN(_0658_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _6115_ (.A1(_0902_),
    .A2(_2897_),
    .B1(_3052_),
    .B2(_2544_),
    .ZN(_0659_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _6116_ (.A1(_0920_),
    .A2(_2897_),
    .B1(_3052_),
    .B2(_2547_),
    .ZN(_0660_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _6117_ (.A1(_0942_),
    .A2(_2897_),
    .B1(_3052_),
    .B2(_2549_),
    .ZN(_0661_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _6118_ (.A1(_0958_),
    .A2(_2897_),
    .B1(_3052_),
    .B2(_2551_),
    .ZN(_0662_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _6119_ (.A1(_0970_),
    .A2(_2897_),
    .B1(_3052_),
    .B2(_2553_),
    .ZN(_0663_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _6120_ (.A1(_0989_),
    .A2(_2897_),
    .B1(_3052_),
    .B2(_2555_),
    .ZN(_0664_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _6121_ (.A1(_1002_),
    .A2(_2897_),
    .B1(_3052_),
    .B2(_2557_),
    .ZN(_0665_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _6122_ (.A1(_1024_),
    .A2(_2896_),
    .B1(_3052_),
    .B2(_2559_),
    .ZN(_0666_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _6123_ (.A1(_1039_),
    .A2(_2896_),
    .B1(_3052_),
    .B2(_2561_),
    .ZN(_0667_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _6124_ (.A1(_1058_),
    .A2(_2896_),
    .B1(_3051_),
    .B2(_2563_),
    .ZN(_0668_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _6125_ (.A1(_1069_),
    .A2(_2896_),
    .B1(_3051_),
    .B2(_2565_),
    .ZN(_0669_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _6126_ (.A1(_1092_),
    .A2(_2896_),
    .B1(_3051_),
    .B2(_2568_),
    .ZN(_0670_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _6127_ (.A1(_1108_),
    .A2(_2896_),
    .B1(_3051_),
    .B2(_2570_),
    .ZN(_0671_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _6128_ (.A1(_1123_),
    .A2(_2896_),
    .B1(_3051_),
    .B2(_2572_),
    .ZN(_0672_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _6129_ (.A1(_1669_),
    .A2(_2896_),
    .B1(_3051_),
    .B2(_2574_),
    .ZN(_0673_));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6130_ (.D(_0010_),
    .CLK(clknet_leaf_8_wb_clk_i),
    .Q(net65));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6131_ (.D(_0011_),
    .CLK(clknet_leaf_8_wb_clk_i),
    .Q(net66));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6132_ (.D(_0012_),
    .CLK(clknet_leaf_1_wb_clk_i),
    .Q(net67));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6133_ (.D(_0013_),
    .CLK(clknet_leaf_2_wb_clk_i),
    .Q(\soc.display_clks_before_active[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6134_ (.D(_0014_),
    .CLK(clknet_4_0_0_wb_clk_i),
    .Q(\soc.video_generator_1.h_count[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _6135_ (.D(_0015_),
    .CLK(clknet_leaf_2_wb_clk_i),
    .Q(\soc.video_generator_1.h_count[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6136_ (.D(_0016_),
    .CLK(clknet_leaf_2_wb_clk_i),
    .Q(\soc.video_generator_1.h_count[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _6137_ (.D(_0017_),
    .CLK(clknet_leaf_1_wb_clk_i),
    .Q(\soc.video_generator_1.h_count[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6138_ (.D(_0018_),
    .CLK(clknet_leaf_1_wb_clk_i),
    .Q(\soc.video_generator_1.h_count[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6139_ (.D(_0019_),
    .CLK(clknet_leaf_1_wb_clk_i),
    .Q(\soc.video_generator_1.h_count[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6140_ (.D(_0020_),
    .CLK(clknet_leaf_1_wb_clk_i),
    .Q(\soc.video_generator_1.h_count[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6141_ (.D(_0021_),
    .CLK(clknet_leaf_0_wb_clk_i),
    .Q(\soc.video_generator_1.h_count[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _6142_ (.D(_0022_),
    .CLK(clknet_leaf_0_wb_clk_i),
    .Q(\soc.video_generator_1.h_count[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6143_ (.D(_0023_),
    .CLK(clknet_leaf_1_wb_clk_i),
    .Q(net64));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6144_ (.D(_0024_),
    .CLK(clknet_leaf_66_wb_clk_i),
    .Q(\soc.ram_encoder_0.output_buffer[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6145_ (.D(_0025_),
    .CLK(clknet_leaf_67_wb_clk_i),
    .Q(\soc.ram_encoder_0.output_buffer[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6146_ (.D(_0026_),
    .CLK(clknet_leaf_67_wb_clk_i),
    .Q(\soc.ram_encoder_0.output_buffer[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6147_ (.D(_0027_),
    .CLK(clknet_leaf_62_wb_clk_i),
    .Q(\soc.ram_encoder_0.output_buffer[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6148_ (.D(_0028_),
    .CLK(clknet_leaf_63_wb_clk_i),
    .Q(\soc.ram_encoder_0.output_buffer[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6149_ (.D(_0029_),
    .CLK(clknet_leaf_62_wb_clk_i),
    .Q(\soc.ram_encoder_0.output_buffer[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6150_ (.D(_0030_),
    .CLK(clknet_leaf_61_wb_clk_i),
    .Q(\soc.ram_encoder_0.output_buffer[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6151_ (.D(_0031_),
    .CLK(clknet_leaf_62_wb_clk_i),
    .Q(\soc.ram_encoder_0.output_buffer[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6152_ (.D(_0032_),
    .CLK(clknet_leaf_61_wb_clk_i),
    .Q(\soc.ram_encoder_0.output_buffer[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6153_ (.D(_0033_),
    .CLK(clknet_leaf_62_wb_clk_i),
    .Q(\soc.ram_encoder_0.output_buffer[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6154_ (.D(_0034_),
    .CLK(clknet_leaf_60_wb_clk_i),
    .Q(\soc.ram_encoder_0.output_buffer[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6155_ (.D(_0035_),
    .CLK(clknet_leaf_44_wb_clk_i),
    .Q(\soc.ram_encoder_0.output_buffer[16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6156_ (.D(_0036_),
    .CLK(clknet_leaf_60_wb_clk_i),
    .Q(\soc.ram_encoder_0.output_buffer[17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6157_ (.D(_0037_),
    .CLK(clknet_leaf_59_wb_clk_i),
    .Q(\soc.ram_encoder_0.output_buffer[18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6158_ (.D(_0038_),
    .CLK(clknet_leaf_60_wb_clk_i),
    .Q(\soc.ram_encoder_0.output_buffer[19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6159_ (.D(_0039_),
    .CLK(clknet_leaf_117_wb_clk_i),
    .Q(\soc.spi_video_ram_1.output_buffer[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6160_ (.D(_0040_),
    .CLK(clknet_leaf_117_wb_clk_i),
    .Q(\soc.spi_video_ram_1.output_buffer[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6161_ (.D(_0041_),
    .CLK(clknet_leaf_117_wb_clk_i),
    .Q(\soc.spi_video_ram_1.output_buffer[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6162_ (.D(_0042_),
    .CLK(clknet_leaf_42_wb_clk_i),
    .Q(\soc.ram_encoder_0.output_bits_left[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6163_ (.D(_0043_),
    .CLK(clknet_leaf_42_wb_clk_i),
    .Q(\soc.ram_encoder_0.output_bits_left[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6164_ (.D(_0044_),
    .CLK(clknet_leaf_44_wb_clk_i),
    .Q(\soc.ram_encoder_0.output_bits_left[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6165_ (.D(_0045_),
    .CLK(clknet_leaf_4_wb_clk_i),
    .Q(\soc.rom_encoder_0.output_bits_left[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6166_ (.D(_0046_),
    .CLK(clknet_leaf_4_wb_clk_i),
    .Q(\soc.rom_encoder_0.output_bits_left[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6167_ (.D(_0047_),
    .CLK(clknet_leaf_4_wb_clk_i),
    .Q(\soc.rom_encoder_0.output_bits_left[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6168_ (.D(_0048_),
    .CLK(net89),
    .Q(\soc.cpu.AReg.data[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6169_ (.D(_0049_),
    .CLK(clknet_leaf_26_wb_clk_i),
    .Q(\soc.rom_encoder_0.output_buffer[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6170_ (.D(_0050_),
    .CLK(clknet_leaf_26_wb_clk_i),
    .Q(\soc.rom_encoder_0.output_buffer[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6171_ (.D(_0051_),
    .CLK(clknet_leaf_26_wb_clk_i),
    .Q(\soc.rom_encoder_0.output_buffer[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6172_ (.D(_0052_),
    .CLK(clknet_leaf_26_wb_clk_i),
    .Q(\soc.rom_encoder_0.output_buffer[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6173_ (.D(_0053_),
    .CLK(clknet_leaf_65_wb_clk_i),
    .Q(\soc.ram_encoder_0.output_buffer[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6174_ (.D(_0054_),
    .CLK(clknet_leaf_67_wb_clk_i),
    .Q(\soc.ram_encoder_0.output_buffer[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6175_ (.D(_0055_),
    .CLK(clknet_leaf_66_wb_clk_i),
    .Q(\soc.ram_encoder_0.output_buffer[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6176_ (.D(_0056_),
    .CLK(clknet_leaf_64_wb_clk_i),
    .Q(\soc.ram_encoder_0.output_buffer[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6177_ (.D(_0057_),
    .CLK(clknet_leaf_134_wb_clk_i),
    .Q(\soc.spi_video_ram_1.output_buffer[23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6178_ (.D(_0058_),
    .CLK(clknet_leaf_114_wb_clk_i),
    .Q(\soc.spi_video_ram_1.output_buffer[22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6179_ (.D(_0059_),
    .CLK(clknet_leaf_134_wb_clk_i),
    .Q(\soc.spi_video_ram_1.output_buffer[21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6180_ (.D(_0060_),
    .CLK(clknet_leaf_134_wb_clk_i),
    .Q(\soc.spi_video_ram_1.output_buffer[20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6181_ (.D(_0061_),
    .CLK(clknet_leaf_134_wb_clk_i),
    .Q(\soc.spi_video_ram_1.output_buffer[19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6182_ (.D(_0062_),
    .CLK(clknet_leaf_114_wb_clk_i),
    .Q(\soc.spi_video_ram_1.output_buffer[18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6183_ (.D(_0063_),
    .CLK(clknet_leaf_113_wb_clk_i),
    .Q(\soc.spi_video_ram_1.output_buffer[17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6184_ (.D(_0064_),
    .CLK(clknet_leaf_113_wb_clk_i),
    .Q(\soc.spi_video_ram_1.output_buffer[16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6185_ (.D(_0065_),
    .CLK(clknet_leaf_135_wb_clk_i),
    .Q(\soc.spi_video_ram_1.output_buffer[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6186_ (.D(_0066_),
    .CLK(clknet_leaf_113_wb_clk_i),
    .Q(\soc.spi_video_ram_1.output_buffer[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6187_ (.D(_0067_),
    .CLK(clknet_leaf_115_wb_clk_i),
    .Q(\soc.spi_video_ram_1.output_buffer[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6188_ (.D(_0068_),
    .CLK(clknet_leaf_110_wb_clk_i),
    .Q(\soc.spi_video_ram_1.output_buffer[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6189_ (.D(_0069_),
    .CLK(clknet_leaf_110_wb_clk_i),
    .Q(\soc.spi_video_ram_1.output_buffer[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6190_ (.D(_0070_),
    .CLK(clknet_leaf_116_wb_clk_i),
    .Q(\soc.spi_video_ram_1.output_buffer[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6191_ (.D(_0071_),
    .CLK(clknet_leaf_116_wb_clk_i),
    .Q(\soc.spi_video_ram_1.output_buffer[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6192_ (.D(_0072_),
    .CLK(clknet_leaf_110_wb_clk_i),
    .Q(\soc.spi_video_ram_1.output_buffer[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6193_ (.D(_0073_),
    .CLK(clknet_leaf_114_wb_clk_i),
    .Q(\soc.spi_video_ram_1.output_buffer[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6194_ (.D(_0074_),
    .CLK(clknet_leaf_113_wb_clk_i),
    .Q(\soc.spi_video_ram_1.output_buffer[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6195_ (.D(_0075_),
    .CLK(clknet_leaf_115_wb_clk_i),
    .Q(\soc.spi_video_ram_1.output_buffer[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6196_ (.D(_0076_),
    .CLK(clknet_leaf_115_wb_clk_i),
    .Q(\soc.spi_video_ram_1.output_buffer[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6197_ (.D(_0077_),
    .CLK(clknet_leaf_133_wb_clk_i),
    .Q(_0000_));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6198_ (.D(_0078_),
    .CLK(clknet_leaf_133_wb_clk_i),
    .Q(_0001_));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6199_ (.D(_0079_),
    .CLK(clknet_leaf_114_wb_clk_i),
    .Q(_0002_));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _6200_ (.D(_0003_),
    .CLK(clknet_leaf_135_wb_clk_i),
    .Q(\soc.spi_video_ram_1.current_state[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6201_ (.D(_0004_),
    .CLK(clknet_leaf_133_wb_clk_i),
    .Q(\soc.spi_video_ram_1.current_state[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _6202_ (.D(_0005_),
    .CLK(clknet_leaf_137_wb_clk_i),
    .Q(\soc.spi_video_ram_1.current_state[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _6203_ (.D(_0006_),
    .CLK(clknet_leaf_135_wb_clk_i),
    .Q(\soc.spi_video_ram_1.current_state[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _6204_ (.D(_0007_),
    .CLK(clknet_leaf_141_wb_clk_i),
    .Q(\soc.spi_video_ram_1.current_state[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6205_ (.D(_0080_),
    .CLK(clknet_leaf_140_wb_clk_i),
    .Q(\soc.spi_video_ram_1.state_counter[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6206_ (.D(_0081_),
    .CLK(clknet_leaf_140_wb_clk_i),
    .Q(\soc.spi_video_ram_1.state_counter[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6207_ (.D(_0082_),
    .CLK(clknet_leaf_139_wb_clk_i),
    .Q(\soc.spi_video_ram_1.state_counter[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6208_ (.D(_0083_),
    .CLK(clknet_leaf_139_wb_clk_i),
    .Q(\soc.spi_video_ram_1.state_counter[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6209_ (.D(_0084_),
    .CLK(clknet_leaf_139_wb_clk_i),
    .Q(\soc.spi_video_ram_1.state_counter[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6210_ (.D(_0085_),
    .CLK(clknet_leaf_139_wb_clk_i),
    .Q(\soc.spi_video_ram_1.state_counter[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6211_ (.D(_0086_),
    .CLK(clknet_leaf_143_wb_clk_i),
    .Q(\soc.spi_video_ram_1.state_counter[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6212_ (.D(_0087_),
    .CLK(clknet_leaf_143_wb_clk_i),
    .Q(\soc.spi_video_ram_1.state_counter[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6213_ (.D(_0088_),
    .CLK(clknet_leaf_140_wb_clk_i),
    .Q(\soc.spi_video_ram_1.state_counter[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6214_ (.D(_0089_),
    .CLK(clknet_leaf_143_wb_clk_i),
    .Q(\soc.spi_video_ram_1.state_counter[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6215_ (.D(_0090_),
    .CLK(clknet_leaf_143_wb_clk_i),
    .Q(\soc.spi_video_ram_1.state_counter[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6216_ (.D(_0091_),
    .CLK(clknet_leaf_9_wb_clk_i),
    .Q(\soc.video_generator_1.v_count[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _6217_ (.D(_0092_),
    .CLK(clknet_leaf_131_wb_clk_i),
    .Q(\soc.video_generator_1.v_count[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _6218_ (.D(_0093_),
    .CLK(clknet_leaf_130_wb_clk_i),
    .Q(\soc.video_generator_1.v_count[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6219_ (.D(_0094_),
    .CLK(clknet_leaf_131_wb_clk_i),
    .Q(\soc.video_generator_1.v_count[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6220_ (.D(_0095_),
    .CLK(clknet_leaf_142_wb_clk_i),
    .Q(\soc.video_generator_1.v_count[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6221_ (.D(_0096_),
    .CLK(clknet_leaf_140_wb_clk_i),
    .Q(\soc.video_generator_1.v_count[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6222_ (.D(_0097_),
    .CLK(clknet_leaf_140_wb_clk_i),
    .Q(\soc.video_generator_1.v_count[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _6223_ (.D(_0098_),
    .CLK(clknet_leaf_142_wb_clk_i),
    .Q(\soc.video_generator_1.v_count[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _6224_ (.D(_0099_),
    .CLK(clknet_leaf_140_wb_clk_i),
    .Q(\soc.video_generator_1.v_count[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6225_ (.D(_0100_),
    .CLK(clknet_leaf_141_wb_clk_i),
    .Q(\soc.video_generator_1.v_count[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _6226_ (.D(_0101_),
    .CLK(clknet_leaf_15_wb_clk_i),
    .Q(\soc.spi_video_ram_1.fifo_in_data[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _6227_ (.D(_0102_),
    .CLK(clknet_leaf_52_wb_clk_i),
    .Q(\soc.spi_video_ram_1.fifo_in_data[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _6228_ (.D(_0103_),
    .CLK(clknet_leaf_16_wb_clk_i),
    .Q(\soc.spi_video_ram_1.fifo_in_data[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _6229_ (.D(_0104_),
    .CLK(clknet_leaf_15_wb_clk_i),
    .Q(\soc.spi_video_ram_1.fifo_in_data[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _6230_ (.D(_0105_),
    .CLK(clknet_leaf_15_wb_clk_i),
    .Q(\soc.spi_video_ram_1.fifo_in_data[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _6231_ (.D(_0106_),
    .CLK(clknet_leaf_52_wb_clk_i),
    .Q(\soc.spi_video_ram_1.fifo_in_data[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _6232_ (.D(_0107_),
    .CLK(clknet_leaf_80_wb_clk_i),
    .Q(\soc.spi_video_ram_1.fifo_in_data[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _6233_ (.D(_0108_),
    .CLK(clknet_leaf_52_wb_clk_i),
    .Q(\soc.spi_video_ram_1.fifo_in_data[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _6234_ (.D(_0109_),
    .CLK(clknet_leaf_80_wb_clk_i),
    .Q(\soc.spi_video_ram_1.fifo_in_data[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _6235_ (.D(_0110_),
    .CLK(clknet_leaf_80_wb_clk_i),
    .Q(\soc.spi_video_ram_1.fifo_in_data[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _6236_ (.D(_0111_),
    .CLK(clknet_leaf_78_wb_clk_i),
    .Q(\soc.spi_video_ram_1.fifo_in_data[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _6237_ (.D(_0112_),
    .CLK(clknet_leaf_74_wb_clk_i),
    .Q(\soc.spi_video_ram_1.fifo_in_data[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _6238_ (.D(_0113_),
    .CLK(clknet_leaf_74_wb_clk_i),
    .Q(\soc.spi_video_ram_1.fifo_in_data[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _6239_ (.D(_0114_),
    .CLK(clknet_leaf_75_wb_clk_i),
    .Q(\soc.spi_video_ram_1.fifo_in_data[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _6240_ (.D(_0115_),
    .CLK(clknet_leaf_78_wb_clk_i),
    .Q(\soc.spi_video_ram_1.fifo_in_data[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _6241_ (.D(_0116_),
    .CLK(clknet_leaf_75_wb_clk_i),
    .Q(\soc.spi_video_ram_1.fifo_in_data[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6242_ (.D(_0117_),
    .CLK(clknet_leaf_12_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[7][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6243_ (.D(_0118_),
    .CLK(clknet_leaf_126_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[7][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6244_ (.D(_0119_),
    .CLK(clknet_leaf_12_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[7][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6245_ (.D(_0120_),
    .CLK(clknet_leaf_14_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[7][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6246_ (.D(_0121_),
    .CLK(clknet_leaf_125_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[7][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6247_ (.D(_0122_),
    .CLK(clknet_leaf_124_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[7][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6248_ (.D(_0123_),
    .CLK(clknet_leaf_122_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[7][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6249_ (.D(_0124_),
    .CLK(clknet_leaf_120_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[7][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6250_ (.D(_0125_),
    .CLK(clknet_leaf_121_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[7][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6251_ (.D(_0126_),
    .CLK(clknet_leaf_81_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[7][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6252_ (.D(_0127_),
    .CLK(clknet_leaf_85_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[7][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6253_ (.D(_0128_),
    .CLK(clknet_leaf_95_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[7][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6254_ (.D(_0129_),
    .CLK(clknet_leaf_91_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[7][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6255_ (.D(_0130_),
    .CLK(clknet_leaf_88_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[7][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6256_ (.D(_0131_),
    .CLK(clknet_leaf_88_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[7][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6257_ (.D(_0132_),
    .CLK(clknet_leaf_93_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[7][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6258_ (.D(_0133_),
    .CLK(clknet_leaf_86_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[7][16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6259_ (.D(_0134_),
    .CLK(clknet_leaf_85_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[7][17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6260_ (.D(_0135_),
    .CLK(clknet_leaf_83_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[7][18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6261_ (.D(_0136_),
    .CLK(clknet_leaf_118_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[7][19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6262_ (.D(_0137_),
    .CLK(clknet_leaf_119_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[7][20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6263_ (.D(_0138_),
    .CLK(clknet_leaf_95_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[7][21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6264_ (.D(_0139_),
    .CLK(clknet_leaf_98_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[7][22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6265_ (.D(_0140_),
    .CLK(clknet_leaf_104_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[7][23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6266_ (.D(_0141_),
    .CLK(clknet_leaf_105_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[7][24] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6267_ (.D(_0142_),
    .CLK(clknet_leaf_111_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[7][25] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6268_ (.D(_0143_),
    .CLK(clknet_leaf_103_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[7][26] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6269_ (.D(_0144_),
    .CLK(clknet_leaf_101_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[7][27] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6270_ (.D(_0145_),
    .CLK(clknet_leaf_117_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[7][28] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6271_ (.D(_0146_),
    .CLK(clknet_leaf_14_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[4][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6272_ (.D(_0147_),
    .CLK(clknet_leaf_128_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[4][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6273_ (.D(_0148_),
    .CLK(clknet_leaf_14_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[4][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6274_ (.D(_0149_),
    .CLK(clknet_leaf_123_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[4][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6275_ (.D(_0150_),
    .CLK(clknet_leaf_124_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[4][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6276_ (.D(_0151_),
    .CLK(clknet_leaf_124_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[4][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6277_ (.D(_0152_),
    .CLK(clknet_leaf_123_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[4][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6278_ (.D(_0153_),
    .CLK(clknet_leaf_125_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[4][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6279_ (.D(_0154_),
    .CLK(clknet_leaf_121_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[4][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6280_ (.D(_0155_),
    .CLK(clknet_leaf_82_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[4][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6281_ (.D(_0156_),
    .CLK(clknet_leaf_90_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[4][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6282_ (.D(_0157_),
    .CLK(clknet_leaf_95_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[4][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6283_ (.D(_0158_),
    .CLK(clknet_leaf_93_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[4][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6284_ (.D(_0159_),
    .CLK(clknet_leaf_87_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[4][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6285_ (.D(_0160_),
    .CLK(clknet_leaf_89_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[4][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6286_ (.D(_0161_),
    .CLK(clknet_leaf_93_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[4][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6287_ (.D(_0162_),
    .CLK(clknet_leaf_121_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[4][16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6288_ (.D(_0163_),
    .CLK(clknet_leaf_85_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[4][17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6289_ (.D(_0164_),
    .CLK(clknet_leaf_82_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[4][18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6290_ (.D(_0165_),
    .CLK(clknet_leaf_87_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[4][19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6291_ (.D(_0166_),
    .CLK(clknet_leaf_119_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[4][20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6292_ (.D(_0167_),
    .CLK(clknet_leaf_96_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[4][21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6293_ (.D(_0168_),
    .CLK(clknet_leaf_89_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[4][22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6294_ (.D(_0169_),
    .CLK(clknet_leaf_104_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[4][23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6295_ (.D(_0170_),
    .CLK(clknet_leaf_106_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[4][24] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6296_ (.D(_0171_),
    .CLK(clknet_leaf_105_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[4][25] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6297_ (.D(_0172_),
    .CLK(clknet_leaf_101_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[4][26] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6298_ (.D(_0173_),
    .CLK(clknet_leaf_97_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[4][27] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6299_ (.D(_0174_),
    .CLK(clknet_leaf_108_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[4][28] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6300_ (.D(_0175_),
    .CLK(clknet_leaf_22_wb_clk_i),
    .Q(\soc.rom_loader.was_loading ));
 gf180mcu_fd_sc_mcu7t5v0__dffnq_2 _6301_ (.D(_0176_),
    .CLKN(clknet_leaf_137_wb_clk_i),
    .Q(\soc.spi_video_ram_1.state_sram_clk_counter[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffnq_2 _6302_ (.D(_0177_),
    .CLKN(clknet_leaf_136_wb_clk_i),
    .Q(\soc.spi_video_ram_1.state_sram_clk_counter[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffnq_1 _6303_ (.D(_0178_),
    .CLKN(clknet_leaf_136_wb_clk_i),
    .Q(\soc.spi_video_ram_1.state_sram_clk_counter[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffnq_1 _6304_ (.D(_0179_),
    .CLKN(clknet_leaf_136_wb_clk_i),
    .Q(\soc.spi_video_ram_1.state_sram_clk_counter[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffnq_1 _6305_ (.D(_0180_),
    .CLKN(clknet_leaf_138_wb_clk_i),
    .Q(\soc.spi_video_ram_1.state_sram_clk_counter[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffnq_1 _6306_ (.D(_0181_),
    .CLKN(clknet_leaf_138_wb_clk_i),
    .Q(\soc.spi_video_ram_1.state_sram_clk_counter[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffnq_1 _6307_ (.D(_0182_),
    .CLKN(clknet_leaf_137_wb_clk_i),
    .Q(\soc.spi_video_ram_1.state_sram_clk_counter[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffnq_2 _6308_ (.D(_0183_),
    .CLKN(clknet_leaf_137_wb_clk_i),
    .Q(\soc.spi_video_ram_1.state_sram_clk_counter[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffnq_2 _6309_ (.D(_0184_),
    .CLKN(clknet_leaf_137_wb_clk_i),
    .Q(\soc.spi_video_ram_1.state_sram_clk_counter[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffnq_1 _6310_ (.D(_0185_),
    .CLKN(clknet_leaf_138_wb_clk_i),
    .Q(net69));
 gf180mcu_fd_sc_mcu7t5v0__dffnq_1 _6311_ (.D(_0186_),
    .CLKN(clknet_leaf_135_wb_clk_i),
    .Q(\soc.spi_video_ram_1.sram_sck_rise_edge ));
 gf180mcu_fd_sc_mcu7t5v0__dffnq_1 _6312_ (.D(_0187_),
    .CLKN(clknet_leaf_140_wb_clk_i),
    .Q(\soc.spi_video_ram_1.sram_sck_fall_edge ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6313_ (.D(_0188_),
    .CLK(clknet_leaf_141_wb_clk_i),
    .Q(net68));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6314_ (.D(_0189_),
    .CLK(clknet_leaf_144_wb_clk_i),
    .Q(\soc.spi_video_ram_1.read_value[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6315_ (.D(_0190_),
    .CLK(clknet_leaf_144_wb_clk_i),
    .Q(\soc.spi_video_ram_1.read_value[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6316_ (.D(_0191_),
    .CLK(clknet_leaf_145_wb_clk_i),
    .Q(\soc.spi_video_ram_1.read_value[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6317_ (.D(_0192_),
    .CLK(clknet_leaf_145_wb_clk_i),
    .Q(\soc.spi_video_ram_1.read_value[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6318_ (.D(_0193_),
    .CLK(clknet_leaf_25_wb_clk_i),
    .Q(\soc.rom_encoder_0.output_buffer[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6319_ (.D(_0194_),
    .CLK(clknet_leaf_25_wb_clk_i),
    .Q(\soc.rom_encoder_0.output_buffer[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6320_ (.D(_0195_),
    .CLK(clknet_leaf_26_wb_clk_i),
    .Q(\soc.rom_encoder_0.output_buffer[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6321_ (.D(_0196_),
    .CLK(clknet_leaf_25_wb_clk_i),
    .Q(\soc.rom_encoder_0.output_buffer[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6322_ (.D(_0197_),
    .CLK(clknet_leaf_25_wb_clk_i),
    .Q(\soc.rom_encoder_0.output_buffer[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6323_ (.D(_0198_),
    .CLK(clknet_leaf_23_wb_clk_i),
    .Q(\soc.rom_encoder_0.output_buffer[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6324_ (.D(_0199_),
    .CLK(clknet_leaf_25_wb_clk_i),
    .Q(\soc.rom_encoder_0.output_buffer[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6325_ (.D(_0200_),
    .CLK(clknet_leaf_24_wb_clk_i),
    .Q(\soc.rom_encoder_0.output_buffer[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6326_ (.D(_0201_),
    .CLK(clknet_leaf_24_wb_clk_i),
    .Q(\soc.rom_encoder_0.output_buffer[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6327_ (.D(_0202_),
    .CLK(clknet_leaf_23_wb_clk_i),
    .Q(\soc.rom_encoder_0.output_buffer[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6328_ (.D(_0203_),
    .CLK(clknet_leaf_23_wb_clk_i),
    .Q(\soc.rom_encoder_0.output_buffer[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6329_ (.D(_0204_),
    .CLK(clknet_leaf_4_wb_clk_i),
    .Q(\soc.rom_encoder_0.output_buffer[16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6330_ (.D(_0205_),
    .CLK(clknet_leaf_24_wb_clk_i),
    .Q(\soc.rom_encoder_0.output_buffer[17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6331_ (.D(_0206_),
    .CLK(clknet_leaf_24_wb_clk_i),
    .Q(\soc.rom_encoder_0.output_buffer[18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6332_ (.D(_0207_),
    .CLK(clknet_leaf_24_wb_clk_i),
    .Q(\soc.rom_encoder_0.output_buffer[19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6333_ (.D(_0208_),
    .CLK(clknet_leaf_112_wb_clk_i),
    .Q(\soc.spi_video_ram_1.buffer_index[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6334_ (.D(_0209_),
    .CLK(clknet_leaf_112_wb_clk_i),
    .Q(\soc.spi_video_ram_1.buffer_index[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6335_ (.D(_0210_),
    .CLK(clknet_leaf_136_wb_clk_i),
    .Q(\soc.spi_video_ram_1.buffer_index[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6336_ (.D(_0211_),
    .CLK(clknet_leaf_136_wb_clk_i),
    .Q(\soc.spi_video_ram_1.buffer_index[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _6337_ (.D(_0212_),
    .CLK(clknet_leaf_112_wb_clk_i),
    .Q(\soc.spi_video_ram_1.buffer_index[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6338_ (.D(_0213_),
    .CLK(clknet_leaf_136_wb_clk_i),
    .Q(\soc.spi_video_ram_1.buffer_index[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6339_ (.D(_0009_),
    .CLK(clknet_leaf_15_wb_clk_i),
    .Q(\soc.spi_video_ram_1.fifo_write_request ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6340_ (.D(_0214_),
    .CLK(clknet_leaf_141_wb_clk_i),
    .Q(\soc.spi_video_ram_1.sram_sio_oe ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _6341_ (.D(_0215_),
    .CLK(clknet_leaf_79_wb_clk_i),
    .Q(\soc.spi_video_ram_1.fifo_in_address[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _6342_ (.D(_0216_),
    .CLK(clknet_leaf_76_wb_clk_i),
    .Q(\soc.spi_video_ram_1.fifo_in_address[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _6343_ (.D(_0217_),
    .CLK(clknet_leaf_78_wb_clk_i),
    .Q(\soc.spi_video_ram_1.fifo_in_address[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _6344_ (.D(_0218_),
    .CLK(clknet_leaf_75_wb_clk_i),
    .Q(\soc.spi_video_ram_1.fifo_in_address[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _6345_ (.D(_0219_),
    .CLK(clknet_leaf_75_wb_clk_i),
    .Q(\soc.spi_video_ram_1.fifo_in_address[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _6346_ (.D(_0220_),
    .CLK(clknet_leaf_76_wb_clk_i),
    .Q(\soc.spi_video_ram_1.fifo_in_address[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _6347_ (.D(_0221_),
    .CLK(clknet_leaf_75_wb_clk_i),
    .Q(\soc.spi_video_ram_1.fifo_in_address[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _6348_ (.D(_0222_),
    .CLK(clknet_4_15_0_wb_clk_i),
    .Q(\soc.spi_video_ram_1.fifo_in_address[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _6349_ (.D(_0223_),
    .CLK(clknet_leaf_76_wb_clk_i),
    .Q(\soc.spi_video_ram_1.fifo_in_address[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _6350_ (.D(_0224_),
    .CLK(clknet_leaf_77_wb_clk_i),
    .Q(\soc.spi_video_ram_1.fifo_in_address[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _6351_ (.D(_0225_),
    .CLK(clknet_leaf_75_wb_clk_i),
    .Q(\soc.spi_video_ram_1.fifo_in_address[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _6352_ (.D(_0226_),
    .CLK(clknet_leaf_76_wb_clk_i),
    .Q(\soc.spi_video_ram_1.fifo_in_address[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _6353_ (.D(_0227_),
    .CLK(clknet_leaf_79_wb_clk_i),
    .Q(\soc.spi_video_ram_1.fifo_in_address[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6354_ (.D(_0008_),
    .CLK(clknet_leaf_133_wb_clk_i),
    .Q(\soc.spi_video_ram_1.fifo_read_request ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6355_ (.D(_0228_),
    .CLK(clknet_leaf_132_wb_clk_i),
    .Q(\soc.spi_video_ram_1.start_read ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6356_ (.D(_0229_),
    .CLK(clknet_leaf_134_wb_clk_i),
    .Q(\soc.spi_video_ram_1.initialized ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6357_ (.D(_0230_),
    .CLK(clknet_leaf_130_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.write_pointer[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6358_ (.D(_0231_),
    .CLK(clknet_leaf_130_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.write_pointer[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _6359_ (.D(_0232_),
    .CLK(clknet_leaf_127_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.write_pointer[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6360_ (.D(_0233_),
    .CLK(clknet_leaf_132_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.read_pointer[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6361_ (.D(_0234_),
    .CLK(clknet_leaf_132_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.read_pointer[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6362_ (.D(_0235_),
    .CLK(clknet_leaf_132_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.read_pointer[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6363_ (.D(_0236_),
    .CLK(clknet_leaf_3_wb_clk_i),
    .Q(\soc.rom_encoder_0.input_bits_left[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6364_ (.D(_0237_),
    .CLK(clknet_leaf_3_wb_clk_i),
    .Q(\soc.rom_encoder_0.input_bits_left[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6365_ (.D(_0238_),
    .CLK(clknet_leaf_3_wb_clk_i),
    .Q(\soc.rom_encoder_0.input_bits_left[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6366_ (.D(_0239_),
    .CLK(clknet_leaf_21_wb_clk_i),
    .Q(\soc.rom_encoder_0.input_buffer[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6367_ (.D(_0240_),
    .CLK(clknet_leaf_21_wb_clk_i),
    .Q(\soc.rom_encoder_0.input_buffer[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6368_ (.D(_0241_),
    .CLK(clknet_leaf_18_wb_clk_i),
    .Q(\soc.rom_encoder_0.input_buffer[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6369_ (.D(_0242_),
    .CLK(clknet_leaf_19_wb_clk_i),
    .Q(\soc.rom_encoder_0.input_buffer[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6370_ (.D(_0243_),
    .CLK(clknet_leaf_18_wb_clk_i),
    .Q(\soc.rom_encoder_0.input_buffer[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6371_ (.D(_0244_),
    .CLK(clknet_leaf_21_wb_clk_i),
    .Q(\soc.rom_encoder_0.input_buffer[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6372_ (.D(_0245_),
    .CLK(clknet_leaf_17_wb_clk_i),
    .Q(\soc.rom_encoder_0.input_buffer[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6373_ (.D(_0246_),
    .CLK(clknet_leaf_16_wb_clk_i),
    .Q(\soc.rom_encoder_0.input_buffer[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6374_ (.D(_0247_),
    .CLK(clknet_leaf_18_wb_clk_i),
    .Q(\soc.rom_encoder_0.input_buffer[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6375_ (.D(_0248_),
    .CLK(clknet_leaf_21_wb_clk_i),
    .Q(\soc.rom_encoder_0.input_buffer[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6376_ (.D(_0249_),
    .CLK(clknet_leaf_17_wb_clk_i),
    .Q(\soc.rom_encoder_0.input_buffer[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6377_ (.D(_0250_),
    .CLK(clknet_leaf_18_wb_clk_i),
    .Q(\soc.rom_encoder_0.input_buffer[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6378_ (.D(_0251_),
    .CLK(clknet_leaf_22_wb_clk_i),
    .Q(\soc.rom_encoder_0.request_write ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6379_ (.D(_0252_),
    .CLK(clknet_leaf_21_wb_clk_i),
    .Q(\soc.rom_encoder_0.request_data_out[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6380_ (.D(_0253_),
    .CLK(clknet_leaf_25_wb_clk_i),
    .Q(\soc.rom_encoder_0.request_data_out[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6381_ (.D(_0254_),
    .CLK(clknet_leaf_11_wb_clk_i),
    .Q(\soc.rom_encoder_0.request_data_out[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6382_ (.D(_0255_),
    .CLK(clknet_leaf_11_wb_clk_i),
    .Q(\soc.rom_encoder_0.request_data_out[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6383_ (.D(_0256_),
    .CLK(clknet_leaf_32_wb_clk_i),
    .Q(\soc.rom_encoder_0.request_data_out[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6384_ (.D(_0257_),
    .CLK(clknet_leaf_32_wb_clk_i),
    .Q(\soc.rom_encoder_0.request_data_out[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6385_ (.D(_0258_),
    .CLK(clknet_leaf_11_wb_clk_i),
    .Q(\soc.rom_encoder_0.request_data_out[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6386_ (.D(_0259_),
    .CLK(clknet_leaf_37_wb_clk_i),
    .Q(\soc.rom_encoder_0.request_data_out[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6387_ (.D(_0260_),
    .CLK(clknet_leaf_11_wb_clk_i),
    .Q(\soc.rom_encoder_0.request_data_out[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6388_ (.D(_0261_),
    .CLK(clknet_leaf_36_wb_clk_i),
    .Q(\soc.rom_encoder_0.request_data_out[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6389_ (.D(_0262_),
    .CLK(clknet_leaf_24_wb_clk_i),
    .Q(\soc.rom_encoder_0.request_data_out[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6390_ (.D(_0263_),
    .CLK(clknet_leaf_37_wb_clk_i),
    .Q(\soc.rom_encoder_0.request_data_out[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6391_ (.D(_0264_),
    .CLK(clknet_leaf_32_wb_clk_i),
    .Q(\soc.rom_encoder_0.request_data_out[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6392_ (.D(_0265_),
    .CLK(clknet_leaf_37_wb_clk_i),
    .Q(\soc.rom_encoder_0.request_data_out[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6393_ (.D(_0266_),
    .CLK(clknet_leaf_11_wb_clk_i),
    .Q(\soc.rom_encoder_0.request_data_out[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6394_ (.D(_0267_),
    .CLK(clknet_leaf_7_wb_clk_i),
    .Q(\soc.rom_encoder_0.request_data_out[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6395_ (.D(_0268_),
    .CLK(clknet_leaf_27_wb_clk_i),
    .Q(\soc.rom_encoder_0.request_address[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6396_ (.D(_0269_),
    .CLK(clknet_leaf_27_wb_clk_i),
    .Q(\soc.rom_encoder_0.request_address[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6397_ (.D(_0270_),
    .CLK(clknet_leaf_27_wb_clk_i),
    .Q(\soc.rom_encoder_0.request_address[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6398_ (.D(_0271_),
    .CLK(clknet_leaf_27_wb_clk_i),
    .Q(\soc.rom_encoder_0.request_address[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6399_ (.D(_0272_),
    .CLK(clknet_leaf_27_wb_clk_i),
    .Q(\soc.rom_encoder_0.request_address[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6400_ (.D(_0273_),
    .CLK(clknet_leaf_32_wb_clk_i),
    .Q(\soc.rom_encoder_0.request_address[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6401_ (.D(_0274_),
    .CLK(clknet_leaf_28_wb_clk_i),
    .Q(\soc.rom_encoder_0.request_address[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6402_ (.D(_0275_),
    .CLK(clknet_leaf_28_wb_clk_i),
    .Q(\soc.rom_encoder_0.request_address[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6403_ (.D(_0276_),
    .CLK(clknet_leaf_20_wb_clk_i),
    .Q(\soc.rom_encoder_0.request_address[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6404_ (.D(_0277_),
    .CLK(clknet_leaf_20_wb_clk_i),
    .Q(\soc.rom_encoder_0.request_address[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6405_ (.D(_0278_),
    .CLK(clknet_leaf_29_wb_clk_i),
    .Q(\soc.rom_encoder_0.request_address[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6406_ (.D(_0279_),
    .CLK(clknet_leaf_21_wb_clk_i),
    .Q(\soc.rom_encoder_0.request_address[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6407_ (.D(_0280_),
    .CLK(clknet_leaf_21_wb_clk_i),
    .Q(\soc.rom_encoder_0.request_address[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6408_ (.D(_0281_),
    .CLK(clknet_leaf_21_wb_clk_i),
    .Q(\soc.rom_encoder_0.request_address[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6409_ (.D(_0282_),
    .CLK(clknet_leaf_23_wb_clk_i),
    .Q(\soc.rom_encoder_0.request_address[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6410_ (.D(_0283_),
    .CLK(clknet_leaf_42_wb_clk_i),
    .Q(net58));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6411_ (.D(_0284_),
    .CLK(clknet_leaf_59_wb_clk_i),
    .Q(net59));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6412_ (.D(_0285_),
    .CLK(clknet_leaf_44_wb_clk_i),
    .Q(net60));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6413_ (.D(_0286_),
    .CLK(clknet_leaf_44_wb_clk_i),
    .Q(net61));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6414_ (.D(_0287_),
    .CLK(clknet_leaf_10_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[3][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6415_ (.D(_0288_),
    .CLK(clknet_leaf_129_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[3][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6416_ (.D(_0289_),
    .CLK(clknet_leaf_10_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[3][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6417_ (.D(_0290_),
    .CLK(clknet_leaf_9_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[3][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6418_ (.D(_0291_),
    .CLK(clknet_leaf_9_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[3][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6419_ (.D(_0292_),
    .CLK(clknet_leaf_129_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[3][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6420_ (.D(_0293_),
    .CLK(clknet_leaf_124_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[3][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6421_ (.D(_0294_),
    .CLK(clknet_leaf_127_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[3][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6422_ (.D(_0295_),
    .CLK(clknet_leaf_114_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[3][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6423_ (.D(_0296_),
    .CLK(clknet_leaf_81_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[3][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6424_ (.D(_0297_),
    .CLK(clknet_leaf_85_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[3][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6425_ (.D(_0298_),
    .CLK(clknet_leaf_92_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[3][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6426_ (.D(_0299_),
    .CLK(clknet_leaf_74_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[3][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6427_ (.D(_0300_),
    .CLK(clknet_leaf_108_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[3][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6428_ (.D(_0301_),
    .CLK(clknet_leaf_99_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[3][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6429_ (.D(_0302_),
    .CLK(clknet_leaf_73_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[3][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6430_ (.D(_0303_),
    .CLK(clknet_leaf_80_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[3][16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6431_ (.D(_0304_),
    .CLK(clknet_leaf_78_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[3][17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6432_ (.D(_0305_),
    .CLK(clknet_leaf_82_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[3][18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6433_ (.D(_0306_),
    .CLK(clknet_leaf_89_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[3][19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6434_ (.D(_0307_),
    .CLK(clknet_leaf_118_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[3][20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6435_ (.D(_0308_),
    .CLK(clknet_leaf_92_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[3][21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6436_ (.D(_0309_),
    .CLK(clknet_leaf_98_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[3][22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6437_ (.D(_0310_),
    .CLK(clknet_leaf_107_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[3][23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6438_ (.D(_0311_),
    .CLK(clknet_leaf_108_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[3][24] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6439_ (.D(_0312_),
    .CLK(clknet_leaf_109_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[3][25] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6440_ (.D(_0313_),
    .CLK(clknet_leaf_100_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[3][26] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6441_ (.D(_0314_),
    .CLK(clknet_leaf_99_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[3][27] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6442_ (.D(_0315_),
    .CLK(clknet_leaf_110_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[3][28] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6443_ (.D(_0316_),
    .CLK(clknet_leaf_7_wb_clk_i),
    .Q(\soc.rom_encoder_0.initialized ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6444_ (.D(_0317_),
    .CLK(clknet_leaf_16_wb_clk_i),
    .Q(\soc.cpu.DMuxJMP.sel[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6445_ (.D(_0318_),
    .CLK(clknet_leaf_51_wb_clk_i),
    .Q(\soc.cpu.DMuxJMP.sel[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6446_ (.D(_0319_),
    .CLK(clknet_leaf_16_wb_clk_i),
    .Q(\soc.cpu.DMuxJMP.sel[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6447_ (.D(_0320_),
    .CLK(clknet_leaf_19_wb_clk_i),
    .Q(\soc.cpu.instruction[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6448_ (.D(_0321_),
    .CLK(clknet_leaf_16_wb_clk_i),
    .Q(\soc.cpu.instruction[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6449_ (.D(_0322_),
    .CLK(clknet_leaf_16_wb_clk_i),
    .Q(\soc.cpu.instruction[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6450_ (.D(_0323_),
    .CLK(clknet_leaf_51_wb_clk_i),
    .Q(\soc.cpu.ALU.no ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6451_ (.D(_0324_),
    .CLK(clknet_leaf_51_wb_clk_i),
    .Q(\soc.cpu.ALU.f ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6452_ (.D(_0325_),
    .CLK(clknet_leaf_51_wb_clk_i),
    .Q(\soc.cpu.ALU.ny ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6453_ (.D(_0326_),
    .CLK(clknet_leaf_51_wb_clk_i),
    .Q(\soc.cpu.ALU.zy ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6454_ (.D(_0327_),
    .CLK(clknet_leaf_51_wb_clk_i),
    .Q(\soc.cpu.ALU.nx ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6455_ (.D(_0328_),
    .CLK(clknet_leaf_16_wb_clk_i),
    .Q(\soc.cpu.ALU.zx ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6456_ (.D(_0329_),
    .CLK(clknet_leaf_48_wb_clk_i),
    .Q(\soc.cpu.instruction[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6457_ (.D(_0330_),
    .CLK(clknet_leaf_19_wb_clk_i),
    .Q(\soc.cpu.instruction[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6458_ (.D(_0331_),
    .CLK(clknet_leaf_16_wb_clk_i),
    .Q(\soc.cpu.instruction[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6459_ (.D(_0332_),
    .CLK(clknet_leaf_19_wb_clk_i),
    .Q(\soc.cpu.instruction[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6460_ (.D(_0333_),
    .CLK(clknet_leaf_7_wb_clk_i),
    .Q(net62));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6461_ (.D(_0334_),
    .CLK(clknet_leaf_7_wb_clk_i),
    .Q(\soc.rom_encoder_0.sram_sio_oe ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6462_ (.D(_0335_),
    .CLK(clknet_leaf_6_wb_clk_i),
    .Q(\soc.rom_encoder_0.current_state[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _6463_ (.D(_0336_),
    .CLK(clknet_leaf_5_wb_clk_i),
    .Q(\soc.rom_encoder_0.current_state[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6464_ (.D(_0337_),
    .CLK(clknet_leaf_5_wb_clk_i),
    .Q(\soc.rom_encoder_0.current_state[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6465_ (.D(_0338_),
    .CLK(clknet_leaf_8_wb_clk_i),
    .Q(\soc.rom_encoder_0.initializing_step[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _6466_ (.D(_0339_),
    .CLK(clknet_leaf_7_wb_clk_i),
    .Q(\soc.rom_encoder_0.initializing_step[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _6467_ (.D(_0340_),
    .CLK(clknet_leaf_3_wb_clk_i),
    .Q(\soc.rom_encoder_0.initializing_step[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _6468_ (.D(_0341_),
    .CLK(clknet_leaf_1_wb_clk_i),
    .Q(\soc.rom_encoder_0.initializing_step[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _6469_ (.D(_0342_),
    .CLK(clknet_leaf_8_wb_clk_i),
    .Q(\soc.rom_encoder_0.initializing_step[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _6470_ (.D(_0343_),
    .CLK(clknet_leaf_35_wb_clk_i),
    .Q(\soc.ram_encoder_0.toggled_sram_sck ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6471_ (.D(_0344_),
    .CLK(clknet_leaf_41_wb_clk_i),
    .Q(\soc.ram_encoder_0.input_bits_left[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6472_ (.D(_0345_),
    .CLK(clknet_leaf_41_wb_clk_i),
    .Q(\soc.ram_encoder_0.input_bits_left[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6473_ (.D(_0346_),
    .CLK(clknet_leaf_41_wb_clk_i),
    .Q(\soc.ram_encoder_0.input_bits_left[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6474_ (.D(_0347_),
    .CLK(clknet_leaf_45_wb_clk_i),
    .Q(\soc.ram_encoder_0.input_buffer[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6475_ (.D(_0348_),
    .CLK(clknet_leaf_58_wb_clk_i),
    .Q(\soc.ram_encoder_0.input_buffer[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6476_ (.D(_0349_),
    .CLK(clknet_leaf_58_wb_clk_i),
    .Q(\soc.ram_encoder_0.input_buffer[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6477_ (.D(_0350_),
    .CLK(clknet_leaf_45_wb_clk_i),
    .Q(\soc.ram_encoder_0.input_buffer[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6478_ (.D(_0351_),
    .CLK(clknet_leaf_45_wb_clk_i),
    .Q(\soc.ram_encoder_0.input_buffer[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6479_ (.D(_0352_),
    .CLK(clknet_leaf_60_wb_clk_i),
    .Q(\soc.ram_encoder_0.input_buffer[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6480_ (.D(_0353_),
    .CLK(clknet_leaf_58_wb_clk_i),
    .Q(\soc.ram_encoder_0.input_buffer[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6481_ (.D(_0354_),
    .CLK(clknet_leaf_46_wb_clk_i),
    .Q(\soc.ram_encoder_0.input_buffer[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6482_ (.D(_0355_),
    .CLK(clknet_leaf_44_wb_clk_i),
    .Q(\soc.ram_encoder_0.input_buffer[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6483_ (.D(_0356_),
    .CLK(clknet_leaf_59_wb_clk_i),
    .Q(\soc.ram_encoder_0.input_buffer[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6484_ (.D(_0357_),
    .CLK(clknet_leaf_59_wb_clk_i),
    .Q(\soc.ram_encoder_0.input_buffer[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6485_ (.D(_0358_),
    .CLK(clknet_leaf_46_wb_clk_i),
    .Q(\soc.ram_encoder_0.input_buffer[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6486_ (.D(_0359_),
    .CLK(clknet_leaf_49_wb_clk_i),
    .Q(\soc.ram_encoder_0.request_write ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6487_ (.D(_0360_),
    .CLK(clknet_leaf_55_wb_clk_i),
    .Q(\soc.ram_encoder_0.request_data_out[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6488_ (.D(_0361_),
    .CLK(clknet_leaf_58_wb_clk_i),
    .Q(\soc.ram_encoder_0.request_data_out[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6489_ (.D(_0362_),
    .CLK(clknet_leaf_63_wb_clk_i),
    .Q(\soc.ram_encoder_0.request_data_out[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6490_ (.D(_0363_),
    .CLK(clknet_leaf_63_wb_clk_i),
    .Q(\soc.ram_encoder_0.request_data_out[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6491_ (.D(_0364_),
    .CLK(clknet_leaf_63_wb_clk_i),
    .Q(\soc.ram_encoder_0.request_data_out[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6492_ (.D(_0365_),
    .CLK(clknet_leaf_61_wb_clk_i),
    .Q(\soc.ram_encoder_0.request_data_out[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6493_ (.D(_0366_),
    .CLK(clknet_leaf_63_wb_clk_i),
    .Q(\soc.ram_encoder_0.request_data_out[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6494_ (.D(_0367_),
    .CLK(clknet_leaf_61_wb_clk_i),
    .Q(\soc.ram_encoder_0.request_data_out[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6495_ (.D(_0368_),
    .CLK(clknet_leaf_43_wb_clk_i),
    .Q(\soc.ram_encoder_0.request_data_out[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6496_ (.D(_0369_),
    .CLK(clknet_leaf_43_wb_clk_i),
    .Q(\soc.ram_encoder_0.request_data_out[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6497_ (.D(_0370_),
    .CLK(clknet_leaf_43_wb_clk_i),
    .Q(\soc.ram_encoder_0.request_data_out[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6498_ (.D(_0371_),
    .CLK(clknet_leaf_46_wb_clk_i),
    .Q(\soc.ram_encoder_0.request_data_out[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6499_ (.D(_0372_),
    .CLK(clknet_leaf_49_wb_clk_i),
    .Q(\soc.ram_encoder_0.request_data_out[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6500_ (.D(_0373_),
    .CLK(clknet_leaf_49_wb_clk_i),
    .Q(\soc.ram_encoder_0.request_data_out[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6501_ (.D(_0374_),
    .CLK(clknet_leaf_49_wb_clk_i),
    .Q(\soc.ram_encoder_0.request_data_out[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6502_ (.D(_0375_),
    .CLK(clknet_leaf_46_wb_clk_i),
    .Q(\soc.ram_encoder_0.request_data_out[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6503_ (.D(_0376_),
    .CLK(clknet_leaf_64_wb_clk_i),
    .Q(\soc.ram_encoder_0.request_address[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6504_ (.D(_0377_),
    .CLK(clknet_leaf_65_wb_clk_i),
    .Q(\soc.ram_encoder_0.request_address[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6505_ (.D(_0378_),
    .CLK(clknet_leaf_64_wb_clk_i),
    .Q(\soc.ram_encoder_0.request_address[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6506_ (.D(_0379_),
    .CLK(clknet_leaf_65_wb_clk_i),
    .Q(\soc.ram_encoder_0.request_address[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6507_ (.D(_0380_),
    .CLK(clknet_leaf_65_wb_clk_i),
    .Q(\soc.ram_encoder_0.request_address[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6508_ (.D(_0381_),
    .CLK(clknet_leaf_66_wb_clk_i),
    .Q(\soc.ram_encoder_0.request_address[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6509_ (.D(_0382_),
    .CLK(clknet_leaf_67_wb_clk_i),
    .Q(\soc.ram_encoder_0.request_address[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6510_ (.D(_0383_),
    .CLK(clknet_leaf_65_wb_clk_i),
    .Q(\soc.ram_encoder_0.request_address[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6511_ (.D(_0384_),
    .CLK(clknet_leaf_65_wb_clk_i),
    .Q(\soc.ram_encoder_0.request_address[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6512_ (.D(_0385_),
    .CLK(clknet_leaf_64_wb_clk_i),
    .Q(\soc.ram_encoder_0.request_address[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6513_ (.D(_0386_),
    .CLK(clknet_4_13_0_wb_clk_i),
    .Q(\soc.ram_encoder_0.request_address[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6514_ (.D(_0387_),
    .CLK(clknet_leaf_66_wb_clk_i),
    .Q(\soc.ram_encoder_0.request_address[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6515_ (.D(_0388_),
    .CLK(clknet_leaf_64_wb_clk_i),
    .Q(\soc.ram_encoder_0.request_address[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6516_ (.D(_0389_),
    .CLK(clknet_leaf_64_wb_clk_i),
    .Q(\soc.ram_encoder_0.request_address[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6517_ (.D(_0390_),
    .CLK(clknet_leaf_60_wb_clk_i),
    .Q(\soc.ram_encoder_0.request_address[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6518_ (.D(_0391_),
    .CLK(clknet_leaf_36_wb_clk_i),
    .Q(\soc.ram_encoder_0.initialized ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6519_ (.D(_0392_),
    .CLK(clknet_leaf_47_wb_clk_i),
    .Q(\soc.ram_data_out[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6520_ (.D(_0393_),
    .CLK(clknet_leaf_47_wb_clk_i),
    .Q(\soc.ram_data_out[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6521_ (.D(_0394_),
    .CLK(clknet_leaf_57_wb_clk_i),
    .Q(\soc.ram_data_out[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6522_ (.D(_0395_),
    .CLK(clknet_leaf_57_wb_clk_i),
    .Q(\soc.ram_data_out[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6523_ (.D(_0396_),
    .CLK(clknet_leaf_56_wb_clk_i),
    .Q(\soc.ram_data_out[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6524_ (.D(_0397_),
    .CLK(clknet_leaf_56_wb_clk_i),
    .Q(\soc.ram_data_out[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6525_ (.D(_0398_),
    .CLK(clknet_leaf_58_wb_clk_i),
    .Q(\soc.ram_data_out[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6526_ (.D(_0399_),
    .CLK(clknet_leaf_55_wb_clk_i),
    .Q(\soc.ram_data_out[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6527_ (.D(_0400_),
    .CLK(clknet_leaf_57_wb_clk_i),
    .Q(\soc.ram_data_out[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6528_ (.D(_0401_),
    .CLK(clknet_leaf_57_wb_clk_i),
    .Q(\soc.ram_data_out[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6529_ (.D(_0402_),
    .CLK(clknet_leaf_57_wb_clk_i),
    .Q(\soc.ram_data_out[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6530_ (.D(_0403_),
    .CLK(clknet_leaf_57_wb_clk_i),
    .Q(\soc.ram_data_out[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6531_ (.D(_0404_),
    .CLK(clknet_leaf_57_wb_clk_i),
    .Q(\soc.ram_data_out[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6532_ (.D(_0405_),
    .CLK(clknet_leaf_47_wb_clk_i),
    .Q(\soc.ram_data_out[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6533_ (.D(_0406_),
    .CLK(clknet_leaf_57_wb_clk_i),
    .Q(\soc.ram_data_out[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6534_ (.D(_0407_),
    .CLK(clknet_leaf_47_wb_clk_i),
    .Q(\soc.ram_data_out[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6535_ (.D(_0408_),
    .CLK(clknet_leaf_39_wb_clk_i),
    .Q(net81));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6536_ (.D(_0409_),
    .CLK(clknet_leaf_40_wb_clk_i),
    .Q(\soc.ram_encoder_0.sram_sio_oe ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6537_ (.D(_0410_),
    .CLK(clknet_leaf_38_wb_clk_i),
    .Q(\soc.ram_encoder_0.current_state[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _6538_ (.D(_0411_),
    .CLK(clknet_leaf_38_wb_clk_i),
    .Q(\soc.ram_encoder_0.current_state[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _6539_ (.D(_0412_),
    .CLK(clknet_leaf_40_wb_clk_i),
    .Q(\soc.ram_encoder_0.current_state[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _6540_ (.D(_0413_),
    .CLK(clknet_leaf_35_wb_clk_i),
    .Q(\soc.ram_encoder_0.initializing_step[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _6541_ (.D(_0414_),
    .CLK(clknet_leaf_34_wb_clk_i),
    .Q(\soc.ram_encoder_0.initializing_step[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _6542_ (.D(_0415_),
    .CLK(clknet_leaf_34_wb_clk_i),
    .Q(\soc.ram_encoder_0.initializing_step[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6543_ (.D(_0416_),
    .CLK(clknet_leaf_34_wb_clk_i),
    .Q(\soc.ram_encoder_0.initializing_step[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6544_ (.D(_0417_),
    .CLK(clknet_leaf_41_wb_clk_i),
    .Q(\soc.ram_encoder_0.initializing_step[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6545_ (.D(_0418_),
    .CLK(clknet_leaf_31_wb_clk_i),
    .Q(\soc.hack_clock_0.counter[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6546_ (.D(_0419_),
    .CLK(clknet_leaf_31_wb_clk_i),
    .Q(\soc.hack_clock_0.counter[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6547_ (.D(_0420_),
    .CLK(clknet_leaf_31_wb_clk_i),
    .Q(\soc.hack_clock_0.counter[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6548_ (.D(_0421_),
    .CLK(clknet_leaf_36_wb_clk_i),
    .Q(\soc.hack_clock_0.counter[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6549_ (.D(_0422_),
    .CLK(clknet_leaf_36_wb_clk_i),
    .Q(\soc.hack_clock_0.counter[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6550_ (.D(_0423_),
    .CLK(clknet_leaf_36_wb_clk_i),
    .Q(\soc.hack_clock_0.counter[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6551_ (.D(_0424_),
    .CLK(clknet_leaf_38_wb_clk_i),
    .Q(\soc.hack_clock_0.counter[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6552_ (.D(_0425_),
    .CLK(clknet_leaf_13_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[5][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6553_ (.D(_0426_),
    .CLK(clknet_leaf_122_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[5][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6554_ (.D(_0427_),
    .CLK(clknet_leaf_17_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[5][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6555_ (.D(_0428_),
    .CLK(clknet_leaf_15_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[5][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6556_ (.D(_0429_),
    .CLK(clknet_leaf_13_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[5][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6557_ (.D(_0430_),
    .CLK(clknet_leaf_122_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[5][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6558_ (.D(_0431_),
    .CLK(clknet_leaf_81_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[5][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6559_ (.D(_0432_),
    .CLK(clknet_leaf_120_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[5][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6560_ (.D(_0433_),
    .CLK(clknet_leaf_121_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[5][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6561_ (.D(_0434_),
    .CLK(clknet_leaf_82_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[5][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6562_ (.D(_0435_),
    .CLK(clknet_leaf_90_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[5][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6563_ (.D(_0436_),
    .CLK(clknet_leaf_94_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[5][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6564_ (.D(_0437_),
    .CLK(clknet_leaf_73_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[5][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6565_ (.D(_0438_),
    .CLK(clknet_leaf_87_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[5][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6566_ (.D(_0439_),
    .CLK(clknet_leaf_85_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[5][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6567_ (.D(_0440_),
    .CLK(clknet_leaf_72_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[5][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6568_ (.D(_0441_),
    .CLK(clknet_leaf_83_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[5][16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6569_ (.D(_0442_),
    .CLK(clknet_leaf_86_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[5][17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6570_ (.D(_0443_),
    .CLK(clknet_leaf_83_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[5][18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6571_ (.D(_0444_),
    .CLK(clknet_leaf_87_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[5][19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6572_ (.D(_0445_),
    .CLK(clknet_leaf_119_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[5][20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6573_ (.D(_0446_),
    .CLK(clknet_leaf_95_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[5][21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6574_ (.D(_0447_),
    .CLK(clknet_leaf_89_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[5][22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6575_ (.D(_0448_),
    .CLK(clknet_leaf_104_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[5][23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6576_ (.D(_0449_),
    .CLK(clknet_leaf_105_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[5][24] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6577_ (.D(_0450_),
    .CLK(clknet_leaf_111_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[5][25] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6578_ (.D(_0451_),
    .CLK(clknet_leaf_103_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[5][26] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6579_ (.D(_0452_),
    .CLK(clknet_4_10_0_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[5][27] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6580_ (.D(_0453_),
    .CLK(clknet_leaf_109_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[5][28] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6581_ (.D(_0454_),
    .CLK(clknet_leaf_11_wb_clk_i),
    .Q(\soc.rom_loader.rom_request ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6582_ (.D(_0455_),
    .CLK(clknet_leaf_6_wb_clk_i),
    .Q(\soc.rom_loader.writing ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6583_ (.D(net20),
    .CLK(clknet_leaf_143_wb_clk_i),
    .Q(\soc.rom_encoder_0.data_out[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6584_ (.D(net21),
    .CLK(clknet_leaf_27_wb_clk_i),
    .Q(\soc.rom_encoder_0.data_out[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6585_ (.D(net22),
    .CLK(clknet_leaf_94_wb_clk_i),
    .Q(\soc.rom_encoder_0.data_out[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6586_ (.D(net23),
    .CLK(clknet_leaf_94_wb_clk_i),
    .Q(\soc.rom_encoder_0.data_out[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6587_ (.D(net24),
    .CLK(clknet_leaf_33_wb_clk_i),
    .Q(\soc.rom_encoder_0.data_out[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6588_ (.D(net25),
    .CLK(clknet_leaf_33_wb_clk_i),
    .Q(\soc.rom_encoder_0.data_out[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6589_ (.D(net26),
    .CLK(clknet_leaf_94_wb_clk_i),
    .Q(\soc.rom_encoder_0.data_out[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6590_ (.D(net27),
    .CLK(clknet_4_13_0_wb_clk_i),
    .Q(\soc.rom_encoder_0.data_out[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6591_ (.D(net28),
    .CLK(clknet_leaf_94_wb_clk_i),
    .Q(\soc.rom_encoder_0.data_out[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6592_ (.D(net30),
    .CLK(clknet_leaf_34_wb_clk_i),
    .Q(\soc.rom_encoder_0.data_out[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6593_ (.D(net31),
    .CLK(clknet_leaf_24_wb_clk_i),
    .Q(\soc.rom_encoder_0.data_out[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6594_ (.D(net32),
    .CLK(clknet_leaf_41_wb_clk_i),
    .Q(\soc.rom_encoder_0.data_out[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6595_ (.D(net33),
    .CLK(clknet_leaf_33_wb_clk_i),
    .Q(\soc.rom_encoder_0.data_out[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6596_ (.D(net34),
    .CLK(clknet_leaf_41_wb_clk_i),
    .Q(\soc.rom_encoder_0.data_out[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6597_ (.D(net35),
    .CLK(clknet_leaf_94_wb_clk_i),
    .Q(\soc.rom_encoder_0.data_out[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6598_ (.D(net36),
    .CLK(clknet_leaf_143_wb_clk_i),
    .Q(\soc.rom_encoder_0.data_out[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6599_ (.D(_0456_),
    .CLK(clknet_leaf_7_wb_clk_i),
    .Q(\soc.rom_encoder_0.toggled_sram_sck ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6600_ (.D(_0457_),
    .CLK(clknet_leaf_29_wb_clk_i),
    .Q(\soc.rom_loader.current_address[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6601_ (.D(_0458_),
    .CLK(clknet_leaf_28_wb_clk_i),
    .Q(\soc.rom_loader.current_address[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6602_ (.D(_0459_),
    .CLK(clknet_leaf_28_wb_clk_i),
    .Q(\soc.rom_loader.current_address[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6603_ (.D(_0460_),
    .CLK(clknet_leaf_28_wb_clk_i),
    .Q(\soc.rom_loader.current_address[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6604_ (.D(_0461_),
    .CLK(clknet_leaf_32_wb_clk_i),
    .Q(\soc.rom_loader.current_address[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6605_ (.D(_0462_),
    .CLK(clknet_leaf_31_wb_clk_i),
    .Q(\soc.rom_loader.current_address[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6606_ (.D(_0463_),
    .CLK(clknet_leaf_31_wb_clk_i),
    .Q(\soc.rom_loader.current_address[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6607_ (.D(_0464_),
    .CLK(clknet_leaf_30_wb_clk_i),
    .Q(\soc.rom_loader.current_address[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6608_ (.D(_0465_),
    .CLK(clknet_leaf_30_wb_clk_i),
    .Q(\soc.rom_loader.current_address[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6609_ (.D(_0466_),
    .CLK(clknet_leaf_29_wb_clk_i),
    .Q(\soc.rom_loader.current_address[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6610_ (.D(_0467_),
    .CLK(clknet_leaf_29_wb_clk_i),
    .Q(\soc.rom_loader.current_address[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6611_ (.D(_0468_),
    .CLK(clknet_leaf_20_wb_clk_i),
    .Q(\soc.rom_loader.current_address[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6612_ (.D(_0469_),
    .CLK(clknet_leaf_20_wb_clk_i),
    .Q(\soc.rom_loader.current_address[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6613_ (.D(_0470_),
    .CLK(clknet_leaf_20_wb_clk_i),
    .Q(\soc.rom_loader.current_address[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6614_ (.D(_0471_),
    .CLK(clknet_leaf_20_wb_clk_i),
    .Q(\soc.rom_loader.current_address[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6615_ (.D(_0472_),
    .CLK(clknet_leaf_6_wb_clk_i),
    .Q(\soc.rom_loader.wait_fall_clk ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6616_ (.D(_0473_),
    .CLK(clknet_leaf_72_wb_clk_i),
    .Q(net83));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _6617_ (.D(\soc.cpu.PC.in[0] ),
    .CLK(net91),
    .Q(\soc.cpu.AReg.data[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _6618_ (.D(\soc.cpu.PC.in[1] ),
    .CLK(net88),
    .Q(\soc.cpu.AReg.data[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6619_ (.D(\soc.cpu.PC.in[2] ),
    .CLK(net87),
    .Q(\soc.cpu.AReg.data[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _6620_ (.D(\soc.cpu.PC.in[3] ),
    .CLK(net87),
    .Q(\soc.cpu.AReg.data[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6621_ (.D(\soc.cpu.PC.in[4] ),
    .CLK(net87),
    .Q(\soc.cpu.AReg.data[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _6622_ (.D(\soc.cpu.PC.in[5] ),
    .CLK(net87),
    .Q(\soc.cpu.AReg.data[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6623_ (.D(\soc.cpu.PC.in[6] ),
    .CLK(net87),
    .Q(\soc.cpu.AReg.data[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6624_ (.D(\soc.cpu.PC.in[7] ),
    .CLK(net88),
    .Q(\soc.cpu.AReg.data[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6625_ (.D(\soc.cpu.PC.in[8] ),
    .CLK(net88),
    .Q(\soc.cpu.AReg.data[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6626_ (.D(\soc.cpu.PC.in[9] ),
    .CLK(net87),
    .Q(\soc.cpu.AReg.data[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _6627_ (.D(\soc.cpu.PC.in[10] ),
    .CLK(net88),
    .Q(\soc.cpu.AReg.data[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _6628_ (.D(\soc.cpu.PC.in[11] ),
    .CLK(net88),
    .Q(\soc.cpu.AReg.data[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _6629_ (.D(\soc.cpu.PC.in[12] ),
    .CLK(net88),
    .Q(\soc.cpu.AReg.data[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _6630_ (.D(\soc.cpu.PC.in[13] ),
    .CLK(net87),
    .Q(\soc.cpu.AReg.data[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _6631_ (.D(\soc.cpu.PC.in[14] ),
    .CLK(net88),
    .Q(\soc.cpu.AReg.data[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6632_ (.D(_0474_),
    .CLK(net89),
    .Q(\soc.cpu.ALU.x[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6633_ (.D(_0475_),
    .CLK(net89),
    .Q(\soc.cpu.ALU.x[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6634_ (.D(_0476_),
    .CLK(net89),
    .Q(\soc.cpu.ALU.x[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6635_ (.D(_0477_),
    .CLK(net89),
    .Q(\soc.cpu.ALU.x[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6636_ (.D(_0478_),
    .CLK(net89),
    .Q(\soc.cpu.ALU.x[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6637_ (.D(_0479_),
    .CLK(net89),
    .Q(\soc.cpu.ALU.x[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6638_ (.D(_0480_),
    .CLK(net89),
    .Q(\soc.cpu.ALU.x[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6639_ (.D(_0481_),
    .CLK(net90),
    .Q(\soc.cpu.ALU.x[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6640_ (.D(_0482_),
    .CLK(net90),
    .Q(\soc.cpu.ALU.x[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6641_ (.D(_0483_),
    .CLK(net90),
    .Q(\soc.cpu.ALU.x[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6642_ (.D(_0484_),
    .CLK(net90),
    .Q(\soc.cpu.ALU.x[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6643_ (.D(_0485_),
    .CLK(net90),
    .Q(\soc.cpu.ALU.x[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6644_ (.D(_0486_),
    .CLK(net90),
    .Q(\soc.cpu.ALU.x[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6645_ (.D(_0487_),
    .CLK(net90),
    .Q(\soc.cpu.ALU.x[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6646_ (.D(_0488_),
    .CLK(net90),
    .Q(\soc.cpu.ALU.x[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6647_ (.D(_0489_),
    .CLK(net89),
    .Q(\soc.cpu.ALU.x[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6648_ (.D(_0490_),
    .CLK(clknet_leaf_12_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[6][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6649_ (.D(_0491_),
    .CLK(clknet_leaf_125_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[6][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6650_ (.D(_0492_),
    .CLK(clknet_leaf_12_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[6][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6651_ (.D(_0493_),
    .CLK(clknet_leaf_15_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[6][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6652_ (.D(_0494_),
    .CLK(clknet_leaf_12_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[6][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6653_ (.D(_0495_),
    .CLK(clknet_leaf_124_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[6][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6654_ (.D(_0496_),
    .CLK(clknet_leaf_123_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[6][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6655_ (.D(_0497_),
    .CLK(clknet_leaf_126_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[6][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6656_ (.D(_0498_),
    .CLK(clknet_leaf_120_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[6][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6657_ (.D(_0499_),
    .CLK(clknet_leaf_80_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[6][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6658_ (.D(_0500_),
    .CLK(clknet_leaf_90_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[6][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6659_ (.D(_0501_),
    .CLK(clknet_leaf_92_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[6][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6660_ (.D(_0502_),
    .CLK(clknet_leaf_91_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[6][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6661_ (.D(_0503_),
    .CLK(clknet_leaf_88_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[6][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6662_ (.D(_0504_),
    .CLK(clknet_leaf_98_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[6][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6663_ (.D(_0505_),
    .CLK(clknet_leaf_93_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[6][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6664_ (.D(_0506_),
    .CLK(clknet_leaf_86_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[6][16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6665_ (.D(_0507_),
    .CLK(clknet_leaf_86_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[6][17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6666_ (.D(_0508_),
    .CLK(clknet_leaf_84_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[6][18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6667_ (.D(_0509_),
    .CLK(clknet_leaf_118_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[6][19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6668_ (.D(_0510_),
    .CLK(clknet_leaf_119_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[6][20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6669_ (.D(_0511_),
    .CLK(clknet_leaf_97_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[6][21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6670_ (.D(_0512_),
    .CLK(clknet_leaf_97_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[6][22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6671_ (.D(_0513_),
    .CLK(clknet_leaf_104_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[6][23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6672_ (.D(_0514_),
    .CLK(clknet_leaf_105_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[6][24] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6673_ (.D(_0515_),
    .CLK(clknet_leaf_111_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[6][25] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6674_ (.D(_0516_),
    .CLK(clknet_leaf_101_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[6][26] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6675_ (.D(_0517_),
    .CLK(clknet_leaf_97_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[6][27] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6676_ (.D(_0518_),
    .CLK(clknet_leaf_116_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[6][28] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6677_ (.D(_0519_),
    .CLK(clknet_leaf_37_wb_clk_i),
    .Q(\soc.cpu.AReg.clk ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6678_ (.D(_0520_),
    .CLK(net84),
    .Q(\soc.cpu.PC.REG.data[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6679_ (.D(_0521_),
    .CLK(net84),
    .Q(\soc.cpu.PC.REG.data[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6680_ (.D(_0522_),
    .CLK(net84),
    .Q(\soc.cpu.PC.REG.data[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6681_ (.D(_0523_),
    .CLK(net84),
    .Q(\soc.cpu.PC.REG.data[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6682_ (.D(_0524_),
    .CLK(net84),
    .Q(\soc.cpu.PC.REG.data[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6683_ (.D(_0525_),
    .CLK(net84),
    .Q(\soc.cpu.PC.REG.data[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6684_ (.D(_0526_),
    .CLK(net85),
    .Q(\soc.cpu.PC.REG.data[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6685_ (.D(_0527_),
    .CLK(net84),
    .Q(\soc.cpu.PC.REG.data[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6686_ (.D(_0528_),
    .CLK(net85),
    .Q(\soc.cpu.PC.REG.data[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6687_ (.D(_0529_),
    .CLK(net85),
    .Q(\soc.cpu.PC.REG.data[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6688_ (.D(_0530_),
    .CLK(net85),
    .Q(\soc.cpu.PC.REG.data[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6689_ (.D(_0531_),
    .CLK(net84),
    .Q(\soc.cpu.PC.REG.data[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6690_ (.D(_0532_),
    .CLK(net86),
    .Q(\soc.cpu.PC.REG.data[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6691_ (.D(_0533_),
    .CLK(net86),
    .Q(\soc.cpu.PC.REG.data[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6692_ (.D(_0534_),
    .CLK(net86),
    .Q(\soc.cpu.PC.REG.data[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6693_ (.D(_0535_),
    .CLK(clknet_leaf_37_wb_clk_i),
    .Q(\soc.hack_clk_strobe ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6694_ (.D(_0536_),
    .CLK(clknet_leaf_50_wb_clk_i),
    .Q(\soc.synch_hack_writeM ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6695_ (.D(_0537_),
    .CLK(clknet_leaf_53_wb_clk_i),
    .Q(\soc.ram_encoder_0.address[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6696_ (.D(_0538_),
    .CLK(clknet_leaf_70_wb_clk_i),
    .Q(\soc.ram_encoder_0.address[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6697_ (.D(_0539_),
    .CLK(clknet_leaf_53_wb_clk_i),
    .Q(\soc.ram_encoder_0.address[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6698_ (.D(_0540_),
    .CLK(clknet_leaf_70_wb_clk_i),
    .Q(\soc.ram_encoder_0.address[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6699_ (.D(_0541_),
    .CLK(clknet_leaf_77_wb_clk_i),
    .Q(\soc.ram_encoder_0.address[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6700_ (.D(_0542_),
    .CLK(clknet_leaf_70_wb_clk_i),
    .Q(\soc.ram_encoder_0.address[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6701_ (.D(_0543_),
    .CLK(clknet_leaf_70_wb_clk_i),
    .Q(\soc.ram_encoder_0.address[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6702_ (.D(_0544_),
    .CLK(clknet_leaf_70_wb_clk_i),
    .Q(\soc.ram_encoder_0.address[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6703_ (.D(_0545_),
    .CLK(clknet_leaf_65_wb_clk_i),
    .Q(\soc.ram_encoder_0.address[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6704_ (.D(_0546_),
    .CLK(clknet_leaf_64_wb_clk_i),
    .Q(\soc.ram_encoder_0.address[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6705_ (.D(_0547_),
    .CLK(clknet_leaf_70_wb_clk_i),
    .Q(\soc.ram_encoder_0.address[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6706_ (.D(_0548_),
    .CLK(clknet_leaf_70_wb_clk_i),
    .Q(\soc.ram_encoder_0.address[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6707_ (.D(_0549_),
    .CLK(clknet_leaf_53_wb_clk_i),
    .Q(\soc.ram_encoder_0.address[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6708_ (.D(_0550_),
    .CLK(clknet_leaf_53_wb_clk_i),
    .Q(\soc.ram_encoder_0.address[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6709_ (.D(_0551_),
    .CLK(clknet_leaf_56_wb_clk_i),
    .Q(\soc.ram_encoder_0.address[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6710_ (.D(_0552_),
    .CLK(clknet_leaf_39_wb_clk_i),
    .Q(\soc.ram_step2_read_request ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6711_ (.D(_0553_),
    .CLK(clknet_leaf_49_wb_clk_i),
    .Q(\soc.ram_step1_write_request ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6712_ (.D(_0554_),
    .CLK(clknet_leaf_6_wb_clk_i),
    .Q(\soc.hack_rom_request ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6713_ (.D(_0555_),
    .CLK(clknet_leaf_8_wb_clk_i),
    .Q(\soc.boot_loading_offset[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _6714_ (.D(_0556_),
    .CLK(clknet_leaf_8_wb_clk_i),
    .Q(\soc.boot_loading_offset[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6715_ (.D(_0557_),
    .CLK(clknet_leaf_9_wb_clk_i),
    .Q(\soc.boot_loading_offset[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _6716_ (.D(_0558_),
    .CLK(clknet_leaf_9_wb_clk_i),
    .Q(\soc.boot_loading_offset[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6717_ (.D(_0559_),
    .CLK(clknet_leaf_8_wb_clk_i),
    .Q(\soc.boot_loading_offset[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6718_ (.D(_0560_),
    .CLK(clknet_leaf_50_wb_clk_i),
    .Q(\soc.rom_encoder_0.write_enable ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6719_ (.D(_0561_),
    .CLK(clknet_leaf_8_wb_clk_i),
    .Q(\soc.hack_wait_clocks[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6720_ (.D(_0562_),
    .CLK(clknet_leaf_8_wb_clk_i),
    .Q(\soc.hack_wait_clocks[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6721_ (.D(_0563_),
    .CLK(net91),
    .Q(net77));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6722_ (.D(_0564_),
    .CLK(net88),
    .Q(net78));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6723_ (.D(_0565_),
    .CLK(net90),
    .Q(net79));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6724_ (.D(_0566_),
    .CLK(net90),
    .Q(net80));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6725_ (.D(_0567_),
    .CLK(net89),
    .Q(\soc.gpio_i_stored[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6726_ (.D(_0568_),
    .CLK(net87),
    .Q(\soc.gpio_i_stored[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6727_ (.D(_0569_),
    .CLK(net91),
    .Q(\soc.gpio_i_stored[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6728_ (.D(_0570_),
    .CLK(net87),
    .Q(\soc.gpio_i_stored[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6729_ (.D(_0571_),
    .CLK(clknet_leaf_10_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[0][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6730_ (.D(_0572_),
    .CLK(clknet_leaf_127_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[0][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6731_ (.D(_0573_),
    .CLK(clknet_leaf_129_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[0][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6732_ (.D(_0574_),
    .CLK(clknet_leaf_129_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[0][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6733_ (.D(_0575_),
    .CLK(clknet_leaf_130_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[0][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6734_ (.D(_0576_),
    .CLK(clknet_leaf_128_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[0][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6735_ (.D(_0577_),
    .CLK(clknet_leaf_124_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[0][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6736_ (.D(_0578_),
    .CLK(clknet_leaf_120_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[0][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6737_ (.D(_0579_),
    .CLK(clknet_leaf_120_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[0][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6738_ (.D(_0580_),
    .CLK(clknet_leaf_122_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[0][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6739_ (.D(_0581_),
    .CLK(clknet_leaf_91_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[0][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6740_ (.D(_0582_),
    .CLK(clknet_leaf_92_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[0][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6741_ (.D(_0583_),
    .CLK(clknet_leaf_73_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[0][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6742_ (.D(_0584_),
    .CLK(clknet_leaf_109_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[0][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6743_ (.D(_0585_),
    .CLK(clknet_leaf_98_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[0][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6744_ (.D(_0586_),
    .CLK(clknet_leaf_73_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[0][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6745_ (.D(_0587_),
    .CLK(clknet_leaf_79_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[0][16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6746_ (.D(_0588_),
    .CLK(clknet_leaf_74_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[0][17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6747_ (.D(_0589_),
    .CLK(clknet_leaf_79_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[0][18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6748_ (.D(_0590_),
    .CLK(clknet_leaf_89_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[0][19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6749_ (.D(_0591_),
    .CLK(clknet_leaf_118_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[0][20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6750_ (.D(_0592_),
    .CLK(clknet_leaf_97_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[0][21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6751_ (.D(_0593_),
    .CLK(clknet_leaf_97_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[0][22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6752_ (.D(_0594_),
    .CLK(clknet_leaf_103_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[0][23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6753_ (.D(_0595_),
    .CLK(clknet_leaf_107_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[0][24] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6754_ (.D(_0596_),
    .CLK(clknet_leaf_107_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[0][25] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6755_ (.D(_0597_),
    .CLK(clknet_leaf_103_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[0][26] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6756_ (.D(_0598_),
    .CLK(clknet_leaf_101_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[0][27] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6757_ (.D(_0599_),
    .CLK(clknet_leaf_110_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[0][28] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6758_ (.D(_0600_),
    .CLK(clknet_leaf_10_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[1][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6759_ (.D(_0601_),
    .CLK(clknet_leaf_126_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[1][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6760_ (.D(_0602_),
    .CLK(clknet_leaf_10_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[1][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6761_ (.D(_0603_),
    .CLK(clknet_leaf_10_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[1][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6762_ (.D(_0604_),
    .CLK(clknet_leaf_130_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[1][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6763_ (.D(_0605_),
    .CLK(clknet_leaf_126_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[1][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6764_ (.D(_0606_),
    .CLK(clknet_leaf_14_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[1][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6765_ (.D(_0607_),
    .CLK(clknet_leaf_127_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[1][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6766_ (.D(_0608_),
    .CLK(clknet_leaf_120_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[1][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6767_ (.D(_0609_),
    .CLK(clknet_leaf_121_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[1][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6768_ (.D(_0610_),
    .CLK(clknet_leaf_85_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[1][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6769_ (.D(_0611_),
    .CLK(clknet_leaf_95_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[1][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6770_ (.D(_0612_),
    .CLK(clknet_leaf_74_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[1][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6771_ (.D(_0613_),
    .CLK(clknet_leaf_88_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[1][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6772_ (.D(_0614_),
    .CLK(clknet_leaf_88_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[1][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6773_ (.D(_0615_),
    .CLK(clknet_leaf_72_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[1][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6774_ (.D(_0616_),
    .CLK(clknet_leaf_79_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[1][16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6775_ (.D(_0617_),
    .CLK(clknet_leaf_74_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[1][17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6776_ (.D(_0618_),
    .CLK(clknet_leaf_84_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[1][18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6777_ (.D(_0619_),
    .CLK(clknet_leaf_89_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[1][19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6778_ (.D(_0620_),
    .CLK(clknet_leaf_88_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[1][20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6779_ (.D(_0621_),
    .CLK(clknet_leaf_96_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[1][21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6780_ (.D(_0622_),
    .CLK(clknet_leaf_97_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[1][22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6781_ (.D(_0623_),
    .CLK(clknet_leaf_104_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[1][23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6782_ (.D(_0624_),
    .CLK(clknet_leaf_107_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[1][24] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6783_ (.D(_0625_),
    .CLK(clknet_leaf_106_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[1][25] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6784_ (.D(_0626_),
    .CLK(clknet_leaf_100_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[1][26] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6785_ (.D(_0627_),
    .CLK(clknet_leaf_98_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[1][27] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6786_ (.D(_0628_),
    .CLK(clknet_leaf_111_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[1][28] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6787_ (.D(_0629_),
    .CLK(clknet_leaf_11_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[2][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6788_ (.D(_0630_),
    .CLK(clknet_leaf_128_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[2][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6789_ (.D(_0631_),
    .CLK(clknet_leaf_10_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[2][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6790_ (.D(_0632_),
    .CLK(clknet_leaf_9_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[2][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6791_ (.D(_0633_),
    .CLK(clknet_leaf_9_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[2][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6792_ (.D(_0634_),
    .CLK(clknet_leaf_128_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[2][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6793_ (.D(_0635_),
    .CLK(clknet_leaf_123_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[2][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6794_ (.D(_0636_),
    .CLK(clknet_leaf_127_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[2][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6795_ (.D(_0637_),
    .CLK(clknet_leaf_115_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[2][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6796_ (.D(_0638_),
    .CLK(clknet_leaf_123_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[2][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6797_ (.D(_0639_),
    .CLK(clknet_leaf_91_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[2][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6798_ (.D(_0640_),
    .CLK(clknet_leaf_90_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[2][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6799_ (.D(_0641_),
    .CLK(clknet_leaf_74_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[2][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6800_ (.D(_0642_),
    .CLK(clknet_leaf_108_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[2][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6801_ (.D(_0643_),
    .CLK(clknet_leaf_99_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[2][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6802_ (.D(_0644_),
    .CLK(clknet_leaf_73_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[2][15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6803_ (.D(_0645_),
    .CLK(clknet_leaf_80_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[2][16] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6804_ (.D(_0646_),
    .CLK(clknet_leaf_84_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[2][17] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6805_ (.D(_0647_),
    .CLK(clknet_leaf_82_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[2][18] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6806_ (.D(_0648_),
    .CLK(clknet_leaf_88_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[2][19] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6807_ (.D(_0649_),
    .CLK(clknet_leaf_119_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[2][20] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6808_ (.D(_0650_),
    .CLK(clknet_leaf_98_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[2][21] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6809_ (.D(_0651_),
    .CLK(clknet_leaf_98_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[2][22] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6810_ (.D(_0652_),
    .CLK(clknet_leaf_106_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[2][23] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6811_ (.D(_0653_),
    .CLK(clknet_leaf_108_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[2][24] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6812_ (.D(_0654_),
    .CLK(clknet_leaf_111_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[2][25] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6813_ (.D(_0655_),
    .CLK(clknet_leaf_99_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[2][26] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6814_ (.D(_0656_),
    .CLK(clknet_leaf_99_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[2][27] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6815_ (.D(_0657_),
    .CLK(clknet_leaf_110_wb_clk_i),
    .Q(\soc.spi_video_ram_1.write_fifo.fifo_mem[2][28] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6816_ (.D(_0658_),
    .CLK(clknet_leaf_55_wb_clk_i),
    .Q(\soc.ram_encoder_0.data_out[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6817_ (.D(_0659_),
    .CLK(clknet_leaf_56_wb_clk_i),
    .Q(\soc.ram_encoder_0.data_out[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6818_ (.D(_0660_),
    .CLK(clknet_leaf_54_wb_clk_i),
    .Q(\soc.ram_encoder_0.data_out[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6819_ (.D(_0661_),
    .CLK(clknet_leaf_54_wb_clk_i),
    .Q(\soc.ram_encoder_0.data_out[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6820_ (.D(_0662_),
    .CLK(clknet_leaf_54_wb_clk_i),
    .Q(\soc.ram_encoder_0.data_out[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6821_ (.D(_0663_),
    .CLK(clknet_leaf_54_wb_clk_i),
    .Q(\soc.ram_encoder_0.data_out[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6822_ (.D(_0664_),
    .CLK(clknet_leaf_54_wb_clk_i),
    .Q(\soc.ram_encoder_0.data_out[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6823_ (.D(_0665_),
    .CLK(clknet_leaf_56_wb_clk_i),
    .Q(\soc.ram_encoder_0.data_out[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6824_ (.D(_0666_),
    .CLK(clknet_leaf_48_wb_clk_i),
    .Q(\soc.ram_encoder_0.data_out[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6825_ (.D(_0667_),
    .CLK(clknet_leaf_48_wb_clk_i),
    .Q(\soc.ram_encoder_0.data_out[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6826_ (.D(_0668_),
    .CLK(clknet_leaf_48_wb_clk_i),
    .Q(\soc.ram_encoder_0.data_out[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6827_ (.D(_0669_),
    .CLK(clknet_leaf_48_wb_clk_i),
    .Q(\soc.ram_encoder_0.data_out[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6828_ (.D(_0670_),
    .CLK(clknet_leaf_50_wb_clk_i),
    .Q(\soc.ram_encoder_0.data_out[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6829_ (.D(_0671_),
    .CLK(clknet_leaf_50_wb_clk_i),
    .Q(\soc.ram_encoder_0.data_out[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6830_ (.D(_0672_),
    .CLK(clknet_leaf_50_wb_clk_i),
    .Q(\soc.ram_encoder_0.data_out[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _6831_ (.D(_0673_),
    .CLK(clknet_leaf_48_wb_clk_i),
    .Q(\soc.ram_encoder_0.data_out[15] ));
 gf180mcu_fd_sc_mcu7t5v0__tieh caravel_hack_soc_226 (.Z(net226));
 gf180mcu_fd_sc_mcu7t5v0__tieh caravel_hack_soc_227 (.Z(net227));
 gf180mcu_fd_sc_mcu7t5v0__tieh caravel_hack_soc_228 (.Z(net228));
 gf180mcu_fd_sc_mcu7t5v0__tieh caravel_hack_soc_229 (.Z(net229));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_0_wb_clk_i (.I(clknet_4_0_0_wb_clk_i),
    .Z(clknet_leaf_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_93 (.ZN(net93));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_94 (.ZN(net94));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_95 (.ZN(net95));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_96 (.ZN(net96));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_97 (.ZN(net97));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_98 (.ZN(net98));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_99 (.ZN(net99));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_100 (.ZN(net100));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_101 (.ZN(net101));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_102 (.ZN(net102));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_103 (.ZN(net103));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_104 (.ZN(net104));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_105 (.ZN(net105));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_106 (.ZN(net106));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_107 (.ZN(net107));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_108 (.ZN(net108));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_109 (.ZN(net109));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_110 (.ZN(net110));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_111 (.ZN(net111));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_112 (.ZN(net112));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_113 (.ZN(net113));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_114 (.ZN(net114));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_115 (.ZN(net115));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_116 (.ZN(net116));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_117 (.ZN(net117));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_118 (.ZN(net118));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_119 (.ZN(net119));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_120 (.ZN(net120));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_121 (.ZN(net121));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_122 (.ZN(net122));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_123 (.ZN(net123));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_124 (.ZN(net124));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_125 (.ZN(net125));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_126 (.ZN(net126));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_127 (.ZN(net127));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_128 (.ZN(net128));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_129 (.ZN(net129));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_130 (.ZN(net130));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_131 (.ZN(net131));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_132 (.ZN(net132));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_133 (.ZN(net133));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_134 (.ZN(net134));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_135 (.ZN(net135));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_136 (.ZN(net136));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_137 (.ZN(net137));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_138 (.ZN(net138));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_139 (.ZN(net139));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_140 (.ZN(net140));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_141 (.ZN(net141));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_142 (.ZN(net142));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_143 (.ZN(net143));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_144 (.ZN(net144));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_145 (.ZN(net145));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_146 (.ZN(net146));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_147 (.ZN(net147));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_148 (.ZN(net148));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_149 (.ZN(net149));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_150 (.ZN(net150));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_151 (.ZN(net151));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_152 (.ZN(net152));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_153 (.ZN(net153));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_154 (.ZN(net154));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_155 (.ZN(net155));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_156 (.ZN(net156));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_157 (.ZN(net157));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_158 (.ZN(net158));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_159 (.ZN(net159));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_160 (.ZN(net160));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_161 (.ZN(net161));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_162 (.ZN(net162));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_163 (.ZN(net163));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_164 (.ZN(net164));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_165 (.ZN(net165));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_166 (.ZN(net166));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_167 (.ZN(net167));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_168 (.ZN(net168));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_169 (.ZN(net169));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_170 (.ZN(net170));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_171 (.ZN(net171));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_172 (.ZN(net172));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_173 (.ZN(net173));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_174 (.ZN(net174));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_175 (.ZN(net175));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_176 (.ZN(net176));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_177 (.ZN(net177));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_178 (.ZN(net178));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_179 (.ZN(net179));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_180 (.ZN(net180));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_181 (.ZN(net181));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_182 (.ZN(net182));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_183 (.ZN(net183));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_184 (.ZN(net184));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_185 (.ZN(net185));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_186 (.ZN(net186));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_187 (.ZN(net187));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_188 (.ZN(net188));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_189 (.ZN(net189));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_190 (.ZN(net190));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_191 (.ZN(net191));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_192 (.ZN(net192));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_193 (.ZN(net193));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_194 (.ZN(net194));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_195 (.ZN(net195));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_196 (.ZN(net196));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_197 (.ZN(net197));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_198 (.ZN(net198));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_199 (.ZN(net199));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_200 (.ZN(net200));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_201 (.ZN(net201));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_202 (.ZN(net202));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_203 (.ZN(net203));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_204 (.ZN(net204));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_205 (.ZN(net205));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_206 (.ZN(net206));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_207 (.ZN(net207));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_208 (.ZN(net208));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_209 (.ZN(net209));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_210 (.ZN(net210));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_211 (.ZN(net211));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_212 (.ZN(net212));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_213 (.ZN(net213));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_214 (.ZN(net214));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_215 (.ZN(net215));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_216 (.ZN(net216));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_217 (.ZN(net217));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_218 (.ZN(net218));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_219 (.ZN(net219));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_220 (.ZN(net220));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_221 (.ZN(net221));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_222 (.ZN(net222));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_223 (.ZN(net223));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_224 (.ZN(net224));
 gf180mcu_fd_sc_mcu7t5v0__tieh caravel_hack_soc_225 (.Z(net225));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6970_ (.I(net49),
    .Z(net46));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6971_ (.I(net49),
    .Z(net47));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6972_ (.I(net49),
    .Z(net48));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6973_ (.I(net53),
    .Z(net50));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6974_ (.I(net53),
    .Z(net51));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6975_ (.I(net53),
    .Z(net52));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6976_ (.I(net57),
    .Z(net54));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6977_ (.I(net57),
    .Z(net55));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6978_ (.I(net57),
    .Z(net56));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_0 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_6 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_7 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_8 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_9 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_10 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_11 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_12 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_13 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_14 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_15 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_16 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_17 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_18 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_19 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_20 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_21 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_22 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_23 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_24 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_25 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_26 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_27 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_28 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_29 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_30 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_31 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_32 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_33 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_34 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_35 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_36 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_37 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_38 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_39 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_40 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_41 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_42 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_43 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_44 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_45 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_46 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_47 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_48 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_49 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_50 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_51 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_52 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_53 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_54 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_55 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_56 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_57 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_58 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_59 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_60 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_61 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_62 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_63 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_64 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_65 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_66 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_67 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_68 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_69 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_70 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_71 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_72 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_73 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_74 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_75 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_76 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_77 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_78 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_79 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_80 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_81 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_82 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_83 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_84 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_85 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_86 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_87 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_88 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_89 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_90 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_91 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_92 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_93 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_94 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_95 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_96 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_97 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_98 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_99 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_100 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_101 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_102 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_103 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_104 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_105 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_106 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_107 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_108 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_109 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_110 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_111 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_112 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_113 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_114 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_115 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_116 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_117 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_118 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_119 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_120 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_121 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_122 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_123 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_124 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_125 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_126 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_127 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_128 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_129 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_130 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_131 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_132 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_133 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_134 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_135 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_136 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_137 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_138 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_139 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_140 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_141 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_142 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_143 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_144 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_145 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_146 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_147 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_148 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_149 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_150 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_151 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_152 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_153 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_154 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_155 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_156 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_157 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_158 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_159 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_160 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_161 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_162 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_163 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_164 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_165 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_166 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_167 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_168 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_169 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_170 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_171 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_172 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_173 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_174 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_175 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_176 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_177 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_178 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_179 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_180 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_181 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_182 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_183 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_184 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_185 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_186 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_187 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_188 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_189 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_190 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_191 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_192 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_193 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_194 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_195 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_196 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_197 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_198 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_199 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_200 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_201 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_202 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_203 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_204 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_205 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_206 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_207 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_208 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_209 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_210 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_211 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_212 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_213 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_214 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_215 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_216 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_217 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_218 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_219 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_220 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_221 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_222 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_223 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_224 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_225 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_226 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_227 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_228 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_229 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_230 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_231 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_232 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_233 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_234 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_235 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_236 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_237 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_238 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_239 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_240 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_241 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_242 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_243 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_244 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_245 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_246 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_247 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_248 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_249 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_250 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_251 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_252 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_253 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_254 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_255 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_256 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_257 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_258 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_259 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_260 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_261 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_262 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_263 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_264 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_265 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_266 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_267 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_268 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_269 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_270 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_271 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_272 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_273 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_274 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_275 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_276 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_277 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_278 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_279 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_280 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_281 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_282 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_283 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_284 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_285 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_286 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_287 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_288 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2420 ();
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 input1 (.I(io_in[10]),
    .Z(net1));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 input2 (.I(io_in[11]),
    .Z(net2));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 input3 (.I(io_in[12]),
    .Z(net3));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 input4 (.I(io_in[13]),
    .Z(net4));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input5 (.I(io_in[16]),
    .Z(net5));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input6 (.I(io_in[17]),
    .Z(net6));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input7 (.I(io_in[18]),
    .Z(net7));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 input8 (.I(io_in[19]),
    .Z(net8));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input9 (.I(io_in[22]),
    .Z(net9));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input10 (.I(io_in[23]),
    .Z(net10));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input11 (.I(io_in[24]),
    .Z(net11));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input12 (.I(io_in[25]),
    .Z(net12));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input13 (.I(io_in[26]),
    .Z(net13));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input14 (.I(io_in[30]),
    .Z(net14));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input15 (.I(io_in[31]),
    .Z(net15));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input16 (.I(io_in[32]),
    .Z(net16));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input17 (.I(io_in[33]),
    .Z(net17));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input18 (.I(la_data_in[0]),
    .Z(net18));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input19 (.I(la_data_in[10]),
    .Z(net19));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input20 (.I(la_data_in[11]),
    .Z(net20));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input21 (.I(la_data_in[12]),
    .Z(net21));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input22 (.I(la_data_in[13]),
    .Z(net22));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input23 (.I(la_data_in[14]),
    .Z(net23));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input24 (.I(la_data_in[15]),
    .Z(net24));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input25 (.I(la_data_in[16]),
    .Z(net25));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input26 (.I(la_data_in[17]),
    .Z(net26));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input27 (.I(la_data_in[18]),
    .Z(net27));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input28 (.I(la_data_in[19]),
    .Z(net28));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input29 (.I(la_data_in[1]),
    .Z(net29));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input30 (.I(la_data_in[20]),
    .Z(net30));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input31 (.I(la_data_in[21]),
    .Z(net31));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input32 (.I(la_data_in[22]),
    .Z(net32));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input33 (.I(la_data_in[23]),
    .Z(net33));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input34 (.I(la_data_in[24]),
    .Z(net34));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input35 (.I(la_data_in[25]),
    .Z(net35));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input36 (.I(la_data_in[26]),
    .Z(net36));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input37 (.I(la_data_in[28]),
    .Z(net37));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input38 (.I(la_data_in[2]),
    .Z(net38));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input39 (.I(la_data_in[3]),
    .Z(net39));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input40 (.I(la_data_in[4]),
    .Z(net40));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input41 (.I(la_data_in[5]),
    .Z(net41));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input42 (.I(la_data_in[6]),
    .Z(net42));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input43 (.I(la_data_in[7]),
    .Z(net43));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input44 (.I(la_data_in[8]),
    .Z(net44));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input45 (.I(la_data_in[9]),
    .Z(net45));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output46 (.I(net46),
    .Z(io_oeb[10]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output47 (.I(net47),
    .Z(io_oeb[11]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output48 (.I(net48),
    .Z(io_oeb[12]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output49 (.I(net49),
    .Z(io_oeb[13]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output50 (.I(net50),
    .Z(io_oeb[16]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output51 (.I(net51),
    .Z(io_oeb[17]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output52 (.I(net52),
    .Z(io_oeb[18]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output53 (.I(net53),
    .Z(io_oeb[19]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output54 (.I(net54),
    .Z(io_oeb[22]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output55 (.I(net55),
    .Z(io_oeb[23]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output56 (.I(net56),
    .Z(io_oeb[24]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output57 (.I(net57),
    .Z(io_oeb[25]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output58 (.I(net58),
    .Z(io_out[10]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output59 (.I(net59),
    .Z(io_out[11]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output60 (.I(net60),
    .Z(io_out[12]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output61 (.I(net61),
    .Z(io_out[13]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output62 (.I(net62),
    .Z(io_out[14]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output63 (.I(net63),
    .Z(io_out[15]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output64 (.I(net64),
    .Z(io_out[16]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output65 (.I(net65),
    .Z(io_out[17]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output66 (.I(net66),
    .Z(io_out[18]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output67 (.I(net67),
    .Z(io_out[19]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output68 (.I(net68),
    .Z(io_out[20]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output69 (.I(net69),
    .Z(io_out[21]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output70 (.I(net70),
    .Z(io_out[22]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output71 (.I(net71),
    .Z(io_out[23]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output72 (.I(net72),
    .Z(io_out[24]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output73 (.I(net73),
    .Z(io_out[25]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output74 (.I(net74),
    .Z(io_out[27]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output75 (.I(net75),
    .Z(io_out[28]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output76 (.I(net76),
    .Z(io_out[29]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output77 (.I(net77),
    .Z(io_out[34]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output78 (.I(net78),
    .Z(io_out[35]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output79 (.I(net79),
    .Z(io_out[36]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output80 (.I(net80),
    .Z(io_out[37]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output81 (.I(net81),
    .Z(io_out[8]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output82 (.I(net82),
    .Z(io_out[9]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output83 (.I(net83),
    .Z(la_data_out[27]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 fanout84 (.I(net86),
    .Z(net84));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 fanout85 (.I(net86),
    .Z(net85));
 gf180mcu_fd_sc_mcu7t5v0__dlyd_1 fanout86 (.I(\soc.cpu.AReg.clk ),
    .Z(net86));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 fanout87 (.I(net88),
    .Z(net87));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 fanout88 (.I(\soc.cpu.AReg.clk ),
    .Z(net88));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 fanout89 (.I(net91),
    .Z(net89));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 fanout90 (.I(net91),
    .Z(net90));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 fanout91 (.I(\soc.cpu.AReg.clk ),
    .Z(net91));
 gf180mcu_fd_sc_mcu7t5v0__tiel caravel_hack_soc_92 (.ZN(net92));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_1_wb_clk_i (.I(clknet_4_0_0_wb_clk_i),
    .Z(clknet_leaf_1_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_2_wb_clk_i (.I(clknet_4_0_0_wb_clk_i),
    .Z(clknet_leaf_2_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_3_wb_clk_i (.I(clknet_4_1_0_wb_clk_i),
    .Z(clknet_leaf_3_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_4_wb_clk_i (.I(clknet_4_1_0_wb_clk_i),
    .Z(clknet_leaf_4_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_5_wb_clk_i (.I(clknet_4_1_0_wb_clk_i),
    .Z(clknet_leaf_5_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_6_wb_clk_i (.I(clknet_4_1_0_wb_clk_i),
    .Z(clknet_leaf_6_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_7_wb_clk_i (.I(clknet_4_1_0_wb_clk_i),
    .Z(clknet_leaf_7_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_8_wb_clk_i (.I(clknet_4_1_0_wb_clk_i),
    .Z(clknet_leaf_8_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_9_wb_clk_i (.I(clknet_4_1_0_wb_clk_i),
    .Z(clknet_leaf_9_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_10_wb_clk_i (.I(clknet_4_1_0_wb_clk_i),
    .Z(clknet_leaf_10_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_11_wb_clk_i (.I(clknet_4_1_0_wb_clk_i),
    .Z(clknet_leaf_11_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_12_wb_clk_i (.I(clknet_4_3_0_wb_clk_i),
    .Z(clknet_leaf_12_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_13_wb_clk_i (.I(clknet_4_3_0_wb_clk_i),
    .Z(clknet_leaf_13_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_14_wb_clk_i (.I(clknet_4_3_0_wb_clk_i),
    .Z(clknet_leaf_14_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_15_wb_clk_i (.I(clknet_4_6_0_wb_clk_i),
    .Z(clknet_leaf_15_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_16_wb_clk_i (.I(clknet_4_6_0_wb_clk_i),
    .Z(clknet_leaf_16_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_17_wb_clk_i (.I(clknet_4_3_0_wb_clk_i),
    .Z(clknet_leaf_17_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_18_wb_clk_i (.I(clknet_4_4_0_wb_clk_i),
    .Z(clknet_leaf_18_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_19_wb_clk_i (.I(clknet_4_4_0_wb_clk_i),
    .Z(clknet_leaf_19_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_20_wb_clk_i (.I(clknet_4_4_0_wb_clk_i),
    .Z(clknet_leaf_20_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_21_wb_clk_i (.I(clknet_4_4_0_wb_clk_i),
    .Z(clknet_leaf_21_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_22_wb_clk_i (.I(clknet_4_4_0_wb_clk_i),
    .Z(clknet_leaf_22_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_23_wb_clk_i (.I(clknet_4_4_0_wb_clk_i),
    .Z(clknet_leaf_23_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_24_wb_clk_i (.I(clknet_4_4_0_wb_clk_i),
    .Z(clknet_leaf_24_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_25_wb_clk_i (.I(clknet_4_5_0_wb_clk_i),
    .Z(clknet_leaf_25_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_26_wb_clk_i (.I(clknet_4_5_0_wb_clk_i),
    .Z(clknet_leaf_26_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_27_wb_clk_i (.I(clknet_4_5_0_wb_clk_i),
    .Z(clknet_leaf_27_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_28_wb_clk_i (.I(clknet_4_5_0_wb_clk_i),
    .Z(clknet_leaf_28_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_29_wb_clk_i (.I(clknet_4_5_0_wb_clk_i),
    .Z(clknet_leaf_29_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_30_wb_clk_i (.I(clknet_4_5_0_wb_clk_i),
    .Z(clknet_leaf_30_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_31_wb_clk_i (.I(clknet_4_5_0_wb_clk_i),
    .Z(clknet_leaf_31_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_32_wb_clk_i (.I(clknet_4_5_0_wb_clk_i),
    .Z(clknet_leaf_32_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_33_wb_clk_i (.I(clknet_4_5_0_wb_clk_i),
    .Z(clknet_leaf_33_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_34_wb_clk_i (.I(clknet_4_7_0_wb_clk_i),
    .Z(clknet_leaf_34_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_35_wb_clk_i (.I(clknet_4_7_0_wb_clk_i),
    .Z(clknet_leaf_35_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_36_wb_clk_i (.I(clknet_4_7_0_wb_clk_i),
    .Z(clknet_leaf_36_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_37_wb_clk_i (.I(clknet_4_7_0_wb_clk_i),
    .Z(clknet_leaf_37_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_38_wb_clk_i (.I(clknet_4_7_0_wb_clk_i),
    .Z(clknet_leaf_38_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_39_wb_clk_i (.I(clknet_4_7_0_wb_clk_i),
    .Z(clknet_leaf_39_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_40_wb_clk_i (.I(clknet_4_7_0_wb_clk_i),
    .Z(clknet_leaf_40_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_41_wb_clk_i (.I(clknet_4_7_0_wb_clk_i),
    .Z(clknet_leaf_41_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_42_wb_clk_i (.I(clknet_4_7_0_wb_clk_i),
    .Z(clknet_leaf_42_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_43_wb_clk_i (.I(clknet_4_7_0_wb_clk_i),
    .Z(clknet_leaf_43_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_44_wb_clk_i (.I(clknet_4_7_0_wb_clk_i),
    .Z(clknet_leaf_44_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_45_wb_clk_i (.I(clknet_4_7_0_wb_clk_i),
    .Z(clknet_leaf_45_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_46_wb_clk_i (.I(clknet_4_6_0_wb_clk_i),
    .Z(clknet_leaf_46_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_47_wb_clk_i (.I(clknet_4_6_0_wb_clk_i),
    .Z(clknet_leaf_47_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_48_wb_clk_i (.I(clknet_4_6_0_wb_clk_i),
    .Z(clknet_leaf_48_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_49_wb_clk_i (.I(clknet_4_6_0_wb_clk_i),
    .Z(clknet_leaf_49_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_50_wb_clk_i (.I(clknet_4_6_0_wb_clk_i),
    .Z(clknet_leaf_50_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_51_wb_clk_i (.I(clknet_4_6_0_wb_clk_i),
    .Z(clknet_leaf_51_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_52_wb_clk_i (.I(clknet_4_6_0_wb_clk_i),
    .Z(clknet_leaf_52_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_53_wb_clk_i (.I(clknet_4_12_0_wb_clk_i),
    .Z(clknet_leaf_53_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_54_wb_clk_i (.I(clknet_4_12_0_wb_clk_i),
    .Z(clknet_leaf_54_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_55_wb_clk_i (.I(clknet_4_13_0_wb_clk_i),
    .Z(clknet_leaf_55_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_56_wb_clk_i (.I(clknet_4_12_0_wb_clk_i),
    .Z(clknet_leaf_56_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_57_wb_clk_i (.I(clknet_4_6_0_wb_clk_i),
    .Z(clknet_leaf_57_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_58_wb_clk_i (.I(clknet_4_13_0_wb_clk_i),
    .Z(clknet_leaf_58_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_59_wb_clk_i (.I(clknet_4_7_0_wb_clk_i),
    .Z(clknet_leaf_59_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_60_wb_clk_i (.I(clknet_4_13_0_wb_clk_i),
    .Z(clknet_leaf_60_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_61_wb_clk_i (.I(clknet_4_13_0_wb_clk_i),
    .Z(clknet_leaf_61_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_62_wb_clk_i (.I(clknet_4_13_0_wb_clk_i),
    .Z(clknet_leaf_62_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_63_wb_clk_i (.I(clknet_4_13_0_wb_clk_i),
    .Z(clknet_leaf_63_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_64_wb_clk_i (.I(clknet_4_12_0_wb_clk_i),
    .Z(clknet_leaf_64_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_65_wb_clk_i (.I(clknet_4_12_0_wb_clk_i),
    .Z(clknet_leaf_65_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_66_wb_clk_i (.I(clknet_4_13_0_wb_clk_i),
    .Z(clknet_leaf_66_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_67_wb_clk_i (.I(clknet_4_13_0_wb_clk_i),
    .Z(clknet_leaf_67_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_70_wb_clk_i (.I(clknet_4_12_0_wb_clk_i),
    .Z(clknet_leaf_70_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_72_wb_clk_i (.I(clknet_4_15_0_wb_clk_i),
    .Z(clknet_leaf_72_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_73_wb_clk_i (.I(clknet_4_15_0_wb_clk_i),
    .Z(clknet_leaf_73_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_74_wb_clk_i (.I(clknet_4_15_0_wb_clk_i),
    .Z(clknet_leaf_74_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_75_wb_clk_i (.I(clknet_4_15_0_wb_clk_i),
    .Z(clknet_leaf_75_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_76_wb_clk_i (.I(clknet_4_15_0_wb_clk_i),
    .Z(clknet_leaf_76_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_77_wb_clk_i (.I(clknet_4_12_0_wb_clk_i),
    .Z(clknet_leaf_77_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_78_wb_clk_i (.I(clknet_4_14_0_wb_clk_i),
    .Z(clknet_leaf_78_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_79_wb_clk_i (.I(clknet_4_14_0_wb_clk_i),
    .Z(clknet_leaf_79_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_80_wb_clk_i (.I(clknet_4_14_0_wb_clk_i),
    .Z(clknet_leaf_80_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_81_wb_clk_i (.I(clknet_4_14_0_wb_clk_i),
    .Z(clknet_leaf_81_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_82_wb_clk_i (.I(clknet_4_9_0_wb_clk_i),
    .Z(clknet_leaf_82_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_83_wb_clk_i (.I(clknet_4_9_0_wb_clk_i),
    .Z(clknet_leaf_83_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_84_wb_clk_i (.I(clknet_4_14_0_wb_clk_i),
    .Z(clknet_leaf_84_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_85_wb_clk_i (.I(clknet_4_9_0_wb_clk_i),
    .Z(clknet_leaf_85_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_86_wb_clk_i (.I(clknet_4_9_0_wb_clk_i),
    .Z(clknet_leaf_86_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_87_wb_clk_i (.I(clknet_4_9_0_wb_clk_i),
    .Z(clknet_leaf_87_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_88_wb_clk_i (.I(clknet_4_9_0_wb_clk_i),
    .Z(clknet_leaf_88_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_89_wb_clk_i (.I(clknet_4_11_0_wb_clk_i),
    .Z(clknet_leaf_89_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_90_wb_clk_i (.I(clknet_4_11_0_wb_clk_i),
    .Z(clknet_leaf_90_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_91_wb_clk_i (.I(clknet_4_14_0_wb_clk_i),
    .Z(clknet_leaf_91_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_92_wb_clk_i (.I(clknet_4_11_0_wb_clk_i),
    .Z(clknet_leaf_92_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_93_wb_clk_i (.I(clknet_4_15_0_wb_clk_i),
    .Z(clknet_leaf_93_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_94_wb_clk_i (.I(clknet_4_11_0_wb_clk_i),
    .Z(clknet_leaf_94_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_95_wb_clk_i (.I(clknet_4_11_0_wb_clk_i),
    .Z(clknet_leaf_95_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_96_wb_clk_i (.I(clknet_4_11_0_wb_clk_i),
    .Z(clknet_leaf_96_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_97_wb_clk_i (.I(clknet_4_11_0_wb_clk_i),
    .Z(clknet_leaf_97_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_98_wb_clk_i (.I(clknet_4_11_0_wb_clk_i),
    .Z(clknet_leaf_98_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_99_wb_clk_i (.I(clknet_4_10_0_wb_clk_i),
    .Z(clknet_leaf_99_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_100_wb_clk_i (.I(clknet_4_10_0_wb_clk_i),
    .Z(clknet_leaf_100_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_101_wb_clk_i (.I(clknet_4_10_0_wb_clk_i),
    .Z(clknet_leaf_101_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_103_wb_clk_i (.I(clknet_4_10_0_wb_clk_i),
    .Z(clknet_leaf_103_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_104_wb_clk_i (.I(clknet_4_10_0_wb_clk_i),
    .Z(clknet_leaf_104_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_105_wb_clk_i (.I(clknet_4_10_0_wb_clk_i),
    .Z(clknet_leaf_105_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_106_wb_clk_i (.I(clknet_4_10_0_wb_clk_i),
    .Z(clknet_leaf_106_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_107_wb_clk_i (.I(clknet_4_10_0_wb_clk_i),
    .Z(clknet_leaf_107_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_108_wb_clk_i (.I(clknet_4_10_0_wb_clk_i),
    .Z(clknet_leaf_108_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_109_wb_clk_i (.I(clknet_4_10_0_wb_clk_i),
    .Z(clknet_leaf_109_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_110_wb_clk_i (.I(clknet_4_8_0_wb_clk_i),
    .Z(clknet_leaf_110_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_111_wb_clk_i (.I(clknet_4_8_0_wb_clk_i),
    .Z(clknet_leaf_111_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_112_wb_clk_i (.I(clknet_4_8_0_wb_clk_i),
    .Z(clknet_leaf_112_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_113_wb_clk_i (.I(clknet_4_8_0_wb_clk_i),
    .Z(clknet_leaf_113_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_114_wb_clk_i (.I(clknet_4_8_0_wb_clk_i),
    .Z(clknet_leaf_114_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_115_wb_clk_i (.I(clknet_4_8_0_wb_clk_i),
    .Z(clknet_leaf_115_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_116_wb_clk_i (.I(clknet_4_8_0_wb_clk_i),
    .Z(clknet_leaf_116_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_117_wb_clk_i (.I(clknet_4_8_0_wb_clk_i),
    .Z(clknet_leaf_117_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_118_wb_clk_i (.I(clknet_4_9_0_wb_clk_i),
    .Z(clknet_leaf_118_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_119_wb_clk_i (.I(clknet_4_9_0_wb_clk_i),
    .Z(clknet_leaf_119_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_120_wb_clk_i (.I(clknet_4_9_0_wb_clk_i),
    .Z(clknet_leaf_120_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_121_wb_clk_i (.I(clknet_4_9_0_wb_clk_i),
    .Z(clknet_leaf_121_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_122_wb_clk_i (.I(clknet_4_9_0_wb_clk_i),
    .Z(clknet_leaf_122_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_123_wb_clk_i (.I(clknet_4_9_0_wb_clk_i),
    .Z(clknet_leaf_123_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_124_wb_clk_i (.I(clknet_4_3_0_wb_clk_i),
    .Z(clknet_leaf_124_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_125_wb_clk_i (.I(clknet_4_3_0_wb_clk_i),
    .Z(clknet_leaf_125_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_126_wb_clk_i (.I(clknet_4_3_0_wb_clk_i),
    .Z(clknet_leaf_126_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_127_wb_clk_i (.I(clknet_4_3_0_wb_clk_i),
    .Z(clknet_leaf_127_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_128_wb_clk_i (.I(clknet_4_3_0_wb_clk_i),
    .Z(clknet_leaf_128_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_129_wb_clk_i (.I(clknet_4_3_0_wb_clk_i),
    .Z(clknet_leaf_129_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_130_wb_clk_i (.I(clknet_4_2_0_wb_clk_i),
    .Z(clknet_leaf_130_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_131_wb_clk_i (.I(clknet_4_2_0_wb_clk_i),
    .Z(clknet_leaf_131_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_132_wb_clk_i (.I(clknet_4_2_0_wb_clk_i),
    .Z(clknet_leaf_132_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_133_wb_clk_i (.I(clknet_4_2_0_wb_clk_i),
    .Z(clknet_leaf_133_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_134_wb_clk_i (.I(clknet_4_2_0_wb_clk_i),
    .Z(clknet_leaf_134_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_135_wb_clk_i (.I(clknet_4_2_0_wb_clk_i),
    .Z(clknet_leaf_135_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_136_wb_clk_i (.I(clknet_4_2_0_wb_clk_i),
    .Z(clknet_leaf_136_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_137_wb_clk_i (.I(clknet_4_2_0_wb_clk_i),
    .Z(clknet_leaf_137_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_138_wb_clk_i (.I(clknet_4_2_0_wb_clk_i),
    .Z(clknet_leaf_138_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_139_wb_clk_i (.I(clknet_4_2_0_wb_clk_i),
    .Z(clknet_leaf_139_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_140_wb_clk_i (.I(clknet_4_2_0_wb_clk_i),
    .Z(clknet_leaf_140_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_141_wb_clk_i (.I(clknet_4_2_0_wb_clk_i),
    .Z(clknet_leaf_141_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_142_wb_clk_i (.I(clknet_4_0_0_wb_clk_i),
    .Z(clknet_leaf_142_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_143_wb_clk_i (.I(clknet_opt_1_0_wb_clk_i),
    .Z(clknet_leaf_143_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_144_wb_clk_i (.I(clknet_4_0_0_wb_clk_i),
    .Z(clknet_leaf_144_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_145_wb_clk_i (.I(clknet_4_0_0_wb_clk_i),
    .Z(clknet_leaf_145_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_0_wb_clk_i (.I(wb_clk_i),
    .Z(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_4_0_0_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_4_0_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_4_1_0_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_4_1_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_4_2_0_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_4_2_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_4_3_0_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_4_3_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_4_4_0_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_4_4_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_4_5_0_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_4_5_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_4_6_0_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_4_6_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_4_7_0_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_4_7_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_4_8_0_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_4_8_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_4_9_0_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_4_9_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_4_10_0_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_4_10_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_4_11_0_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_4_11_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_4_12_0_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_4_12_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_4_13_0_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_4_13_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_4_14_0_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_4_14_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_4_15_0_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_4_15_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_opt_1_0_wb_clk_i (.I(clknet_4_0_0_wb_clk_i),
    .Z(clknet_opt_1_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_1 (.I(net22));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_2 (.I(net25));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_3 (.I(net72));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_4 (.I(net81));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_13 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_1_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_1_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_1_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_1_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_1_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_1_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_3_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_4_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_4_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_5_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_5_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_5_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_5_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_5_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_6_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_6_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_6_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_7_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_7_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_7_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_7_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_7_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_8_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_8_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_8_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_9_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_9_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_15 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_10_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_10_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_10_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_11_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_11_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_11_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_12_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_12_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_13_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_13_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_13_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_14_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_14_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_14_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_14_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_14_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_14_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_14_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_14_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_14_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_15_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_15_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_15_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_16_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_16_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_17_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_17_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_17_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_17_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_17_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_17_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_17_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_17_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_17_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_18_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_18_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_18_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_18_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_18_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_19_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_19_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_19_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_19_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_20_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_20_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_20_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_20_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_20_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_20_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_20_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_21_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_21_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_21_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_22_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_22_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_22_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_23_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_23_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_24_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_24_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_24_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_24_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_24_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_24_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_24_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_25_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_25_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_25_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_25_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_25_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_26_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_26_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_27_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_27_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_27_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_27_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_28_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_28_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_28_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_28_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_29_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_29_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_29_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_30_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_30_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_30_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_30_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_31_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_32_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_32_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_32_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_32_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_33_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_34_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_34_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_34_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_36_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_36_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_36_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_37_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_38_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_39_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_39_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_39_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_39_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_40_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_40_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_40_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_40_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_40_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_40_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_40_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_41_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_43_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_45_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_45_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_45_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_45_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_45_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_47_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_47_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_48_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_49_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_50_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_51_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_55_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_56_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_59_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_62_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_62_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_62_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_64_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_65_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_66_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_66_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_67_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_67_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_68_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_69_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_69_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_69_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_70_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_70_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_71_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_72_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_72_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_72_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_73_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_73_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_75_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_76_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_76_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_76_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_76_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_76_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_77_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_77_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_77_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_78_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_78_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_78_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_79_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_79_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_80_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_80_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_80_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_80_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_81_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_81_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_81_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_82_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_82_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_83_15 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_83_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_83_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_84_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_84_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_85_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_85_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_85_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_85_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_86_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_87_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_87_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_87_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_88_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_88_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_88_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_89_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_89_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_89_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_90_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_90_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_90_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_91_15 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_91_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_91_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_92_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_93_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_93_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_93_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_94_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_94_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_94_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_94_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_95_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_96_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_96_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_96_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_96_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_97_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_97_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_98_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_99_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_99_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_15 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_100_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_100_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_101_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_101_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_101_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_102_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_103_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_103_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_103_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_104_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_104_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_105_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_105_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_106_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_106_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_107_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_107_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_107_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_108_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_108_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_109_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_109_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_109_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_15 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_110_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_110_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_111_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_111_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_112_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_112_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_112_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_113_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_114_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_114_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_115_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_15 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_116_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_116_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_116_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_117_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_117_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_118_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_118_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_119_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_119_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_120_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_120_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_121_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_121_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_122_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_122_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_122_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_123_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_123_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_124_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_124_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_124_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_126_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_126_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_127_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_127_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_128_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_129_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_132_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_133_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_134_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_135_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_135_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_136_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_137_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_138_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_138_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_138_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_139_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_139_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_140_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_141_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_141_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_142_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_142_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_142_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_142_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_142_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_143_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_143_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_143_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_143_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_143_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_143_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_143_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_143_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_143_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_144_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1043 ();
 assign io_oeb[0] = net92;
 assign io_oeb[14] = net102;
 assign io_oeb[15] = net103;
 assign io_oeb[1] = net93;
 assign io_oeb[20] = net104;
 assign io_oeb[21] = net105;
 assign io_oeb[26] = net225;
 assign io_oeb[27] = net106;
 assign io_oeb[28] = net107;
 assign io_oeb[29] = net108;
 assign io_oeb[2] = net94;
 assign io_oeb[30] = net226;
 assign io_oeb[31] = net227;
 assign io_oeb[32] = net228;
 assign io_oeb[33] = net229;
 assign io_oeb[34] = net109;
 assign io_oeb[35] = net110;
 assign io_oeb[36] = net111;
 assign io_oeb[37] = net112;
 assign io_oeb[3] = net95;
 assign io_oeb[4] = net96;
 assign io_oeb[5] = net97;
 assign io_oeb[6] = net98;
 assign io_oeb[7] = net99;
 assign io_oeb[8] = net100;
 assign io_oeb[9] = net101;
 assign io_out[0] = net113;
 assign io_out[1] = net114;
 assign io_out[26] = net121;
 assign io_out[2] = net115;
 assign io_out[30] = net122;
 assign io_out[31] = net123;
 assign io_out[32] = net124;
 assign io_out[33] = net125;
 assign io_out[3] = net116;
 assign io_out[4] = net117;
 assign io_out[5] = net118;
 assign io_out[6] = net119;
 assign io_out[7] = net120;
 assign irq[0] = net126;
 assign irq[1] = net127;
 assign irq[2] = net128;
 assign la_data_out[0] = net129;
 assign la_data_out[10] = net139;
 assign la_data_out[11] = net140;
 assign la_data_out[12] = net141;
 assign la_data_out[13] = net142;
 assign la_data_out[14] = net143;
 assign la_data_out[15] = net144;
 assign la_data_out[16] = net145;
 assign la_data_out[17] = net146;
 assign la_data_out[18] = net147;
 assign la_data_out[19] = net148;
 assign la_data_out[1] = net130;
 assign la_data_out[20] = net149;
 assign la_data_out[21] = net150;
 assign la_data_out[22] = net151;
 assign la_data_out[23] = net152;
 assign la_data_out[24] = net153;
 assign la_data_out[25] = net154;
 assign la_data_out[26] = net155;
 assign la_data_out[28] = net156;
 assign la_data_out[29] = net157;
 assign la_data_out[2] = net131;
 assign la_data_out[30] = net158;
 assign la_data_out[31] = net159;
 assign la_data_out[32] = net160;
 assign la_data_out[33] = net161;
 assign la_data_out[34] = net162;
 assign la_data_out[35] = net163;
 assign la_data_out[36] = net164;
 assign la_data_out[37] = net165;
 assign la_data_out[38] = net166;
 assign la_data_out[39] = net167;
 assign la_data_out[3] = net132;
 assign la_data_out[40] = net168;
 assign la_data_out[41] = net169;
 assign la_data_out[42] = net170;
 assign la_data_out[43] = net171;
 assign la_data_out[44] = net172;
 assign la_data_out[45] = net173;
 assign la_data_out[46] = net174;
 assign la_data_out[47] = net175;
 assign la_data_out[48] = net176;
 assign la_data_out[49] = net177;
 assign la_data_out[4] = net133;
 assign la_data_out[50] = net178;
 assign la_data_out[51] = net179;
 assign la_data_out[52] = net180;
 assign la_data_out[53] = net181;
 assign la_data_out[54] = net182;
 assign la_data_out[55] = net183;
 assign la_data_out[56] = net184;
 assign la_data_out[57] = net185;
 assign la_data_out[58] = net186;
 assign la_data_out[59] = net187;
 assign la_data_out[5] = net134;
 assign la_data_out[60] = net188;
 assign la_data_out[61] = net189;
 assign la_data_out[62] = net190;
 assign la_data_out[63] = net191;
 assign la_data_out[6] = net135;
 assign la_data_out[7] = net136;
 assign la_data_out[8] = net137;
 assign la_data_out[9] = net138;
 assign wbs_ack_o = net192;
 assign wbs_dat_o[0] = net193;
 assign wbs_dat_o[10] = net203;
 assign wbs_dat_o[11] = net204;
 assign wbs_dat_o[12] = net205;
 assign wbs_dat_o[13] = net206;
 assign wbs_dat_o[14] = net207;
 assign wbs_dat_o[15] = net208;
 assign wbs_dat_o[16] = net209;
 assign wbs_dat_o[17] = net210;
 assign wbs_dat_o[18] = net211;
 assign wbs_dat_o[19] = net212;
 assign wbs_dat_o[1] = net194;
 assign wbs_dat_o[20] = net213;
 assign wbs_dat_o[21] = net214;
 assign wbs_dat_o[22] = net215;
 assign wbs_dat_o[23] = net216;
 assign wbs_dat_o[24] = net217;
 assign wbs_dat_o[25] = net218;
 assign wbs_dat_o[26] = net219;
 assign wbs_dat_o[27] = net220;
 assign wbs_dat_o[28] = net221;
 assign wbs_dat_o[29] = net222;
 assign wbs_dat_o[2] = net195;
 assign wbs_dat_o[30] = net223;
 assign wbs_dat_o[31] = net224;
 assign wbs_dat_o[3] = net196;
 assign wbs_dat_o[4] = net197;
 assign wbs_dat_o[5] = net198;
 assign wbs_dat_o[6] = net199;
 assign wbs_dat_o[7] = net200;
 assign wbs_dat_o[8] = net201;
 assign wbs_dat_o[9] = net202;
endmodule

