* NGSPICE file created from caravel_hack_soc.ext - technology: gf180mcuC

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_4 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_1 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_1 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_16 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_1 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffq_1 D CLK Q VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__tieh abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__tieh Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__tiel abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__tiel ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux2_2 I0 I1 S Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_32 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_32 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_2 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__filltie abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__filltie VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_8 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_64 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_64 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai32_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai32_1 A1 A2 A3 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffq_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffq_2 D CLK Q VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_1 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_2 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux4_1 I0 I1 I2 I3 S0 S1 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_2 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_2 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_4 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_1 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_1 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_1 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and3_1 A1 A2 A3 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_1 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_1 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_1 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_3 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_3 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_1 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_1 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and4_1 A1 A2 A3 A4 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_4 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xnor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xnor2_1 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffnq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffnq_1 D CLKN Q VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai31_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_1 A1 A2 A3 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__endcap abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__endcap VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_1 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_4 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_1 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor2_1 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_2 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and2_1 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_2 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai31_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_2 A1 A2 A3 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or2_1 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_4 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_1 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai22_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_1 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_4 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and3_2 A1 A2 A3 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_2 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_2 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or3_2 A1 A2 A3 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_3 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_3 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or4_1 A1 A2 A3 A4 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai221_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai221_1 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_2 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_4 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_4 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_2 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_4 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor3_1 A1 A2 A3 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xnor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xnor3_1 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_2 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or3_1 A1 A2 A3 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xnor2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xnor2_2 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dlyd_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dlyd_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_2 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_2 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_4 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai221_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai221_2 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dlyc_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dlyc_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffnq_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffnq_2 D CLKN Q VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai32_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai32_2 A1 A2 A3 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_4 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor3_2 A1 A2 A3 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffq_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffq_4 D CLK Q VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dlyb_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dlyb_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_4 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi222_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi222_1 A1 A2 B1 B2 C1 C2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xnor3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xnor3_2 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai31_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_4 A1 A2 A3 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and2_2 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai222_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai222_2 A1 A2 B1 B2 C1 C2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_4 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor2_2 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_2 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_2 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and4_2 A1 A2 A3 A4 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__antenna abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__antenna I VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_3 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_3 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai22_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_2 A1 A2 B1 B2 ZN VDD VSS
.ends

.subckt caravel_hack_soc io_in[0] io_in[10] io_in[11] io_in[12] io_in[13] io_in[14]
+ io_in[15] io_in[16] io_in[17] io_in[18] io_in[19] io_in[1] io_in[20] io_in[21] io_in[22]
+ io_in[23] io_in[24] io_in[25] io_in[26] io_in[27] io_in[28] io_in[29] io_in[2] io_in[30]
+ io_in[31] io_in[32] io_in[33] io_in[34] io_in[35] io_in[36] io_in[37] io_in[3] io_in[4]
+ io_in[5] io_in[6] io_in[7] io_in[8] io_in[9] io_oeb[0] io_oeb[10] io_oeb[11] io_oeb[12]
+ io_oeb[13] io_oeb[14] io_oeb[15] io_oeb[16] io_oeb[17] io_oeb[18] io_oeb[19] io_oeb[1]
+ io_oeb[20] io_oeb[21] io_oeb[22] io_oeb[23] io_oeb[24] io_oeb[25] io_oeb[26] io_oeb[27]
+ io_oeb[28] io_oeb[29] io_oeb[2] io_oeb[30] io_oeb[31] io_oeb[32] io_oeb[33] io_oeb[34]
+ io_oeb[35] io_oeb[36] io_oeb[37] io_oeb[3] io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7]
+ io_oeb[8] io_oeb[9] io_out[0] io_out[10] io_out[11] io_out[12] io_out[13] io_out[14]
+ io_out[15] io_out[16] io_out[17] io_out[18] io_out[19] io_out[1] io_out[20] io_out[21]
+ io_out[22] io_out[23] io_out[24] io_out[25] io_out[26] io_out[27] io_out[28] io_out[29]
+ io_out[2] io_out[30] io_out[31] io_out[32] io_out[33] io_out[34] io_out[35] io_out[36]
+ io_out[37] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7] io_out[8] io_out[9]
+ irq[0] irq[1] irq[2] la_data_in[0] la_data_in[10] la_data_in[11] la_data_in[12]
+ la_data_in[13] la_data_in[14] la_data_in[15] la_data_in[16] la_data_in[17] la_data_in[18]
+ la_data_in[19] la_data_in[1] la_data_in[20] la_data_in[21] la_data_in[22] la_data_in[23]
+ la_data_in[24] la_data_in[25] la_data_in[26] la_data_in[27] la_data_in[28] la_data_in[29]
+ la_data_in[2] la_data_in[30] la_data_in[31] la_data_in[32] la_data_in[33] la_data_in[34]
+ la_data_in[35] la_data_in[36] la_data_in[37] la_data_in[38] la_data_in[39] la_data_in[3]
+ la_data_in[40] la_data_in[41] la_data_in[42] la_data_in[43] la_data_in[44] la_data_in[45]
+ la_data_in[46] la_data_in[47] la_data_in[48] la_data_in[49] la_data_in[4] la_data_in[50]
+ la_data_in[51] la_data_in[52] la_data_in[53] la_data_in[54] la_data_in[55] la_data_in[56]
+ la_data_in[57] la_data_in[58] la_data_in[59] la_data_in[5] la_data_in[60] la_data_in[61]
+ la_data_in[62] la_data_in[63] la_data_in[6] la_data_in[7] la_data_in[8] la_data_in[9]
+ la_data_out[0] la_data_out[10] la_data_out[11] la_data_out[12] la_data_out[13] la_data_out[14]
+ la_data_out[15] la_data_out[16] la_data_out[17] la_data_out[18] la_data_out[19]
+ la_data_out[1] la_data_out[20] la_data_out[21] la_data_out[22] la_data_out[23] la_data_out[24]
+ la_data_out[25] la_data_out[26] la_data_out[27] la_data_out[28] la_data_out[29]
+ la_data_out[2] la_data_out[30] la_data_out[31] la_data_out[32] la_data_out[33] la_data_out[34]
+ la_data_out[35] la_data_out[36] la_data_out[37] la_data_out[38] la_data_out[39]
+ la_data_out[3] la_data_out[40] la_data_out[41] la_data_out[42] la_data_out[43] la_data_out[44]
+ la_data_out[45] la_data_out[46] la_data_out[47] la_data_out[48] la_data_out[49]
+ la_data_out[4] la_data_out[50] la_data_out[51] la_data_out[52] la_data_out[53] la_data_out[54]
+ la_data_out[55] la_data_out[56] la_data_out[57] la_data_out[58] la_data_out[59]
+ la_data_out[5] la_data_out[60] la_data_out[61] la_data_out[62] la_data_out[63] la_data_out[6]
+ la_data_out[7] la_data_out[8] la_data_out[9] la_oenb[0] la_oenb[10] la_oenb[11]
+ la_oenb[12] la_oenb[13] la_oenb[14] la_oenb[15] la_oenb[16] la_oenb[17] la_oenb[18]
+ la_oenb[19] la_oenb[1] la_oenb[20] la_oenb[21] la_oenb[22] la_oenb[23] la_oenb[24]
+ la_oenb[25] la_oenb[26] la_oenb[27] la_oenb[28] la_oenb[29] la_oenb[2] la_oenb[30]
+ la_oenb[31] la_oenb[32] la_oenb[33] la_oenb[34] la_oenb[35] la_oenb[36] la_oenb[37]
+ la_oenb[38] la_oenb[39] la_oenb[3] la_oenb[40] la_oenb[41] la_oenb[42] la_oenb[43]
+ la_oenb[44] la_oenb[45] la_oenb[46] la_oenb[47] la_oenb[48] la_oenb[49] la_oenb[4]
+ la_oenb[50] la_oenb[51] la_oenb[52] la_oenb[53] la_oenb[54] la_oenb[55] la_oenb[56]
+ la_oenb[57] la_oenb[58] la_oenb[59] la_oenb[5] la_oenb[60] la_oenb[61] la_oenb[62]
+ la_oenb[63] la_oenb[6] la_oenb[7] la_oenb[8] la_oenb[9] vdd vss wb_clk_i wb_rst_i
+ wbs_ack_o wbs_adr_i[0] wbs_adr_i[10] wbs_adr_i[11] wbs_adr_i[12] wbs_adr_i[13] wbs_adr_i[14]
+ wbs_adr_i[15] wbs_adr_i[16] wbs_adr_i[17] wbs_adr_i[18] wbs_adr_i[19] wbs_adr_i[1]
+ wbs_adr_i[20] wbs_adr_i[21] wbs_adr_i[22] wbs_adr_i[23] wbs_adr_i[24] wbs_adr_i[25]
+ wbs_adr_i[26] wbs_adr_i[27] wbs_adr_i[28] wbs_adr_i[29] wbs_adr_i[2] wbs_adr_i[30]
+ wbs_adr_i[31] wbs_adr_i[3] wbs_adr_i[4] wbs_adr_i[5] wbs_adr_i[6] wbs_adr_i[7] wbs_adr_i[8]
+ wbs_adr_i[9] wbs_cyc_i wbs_dat_i[0] wbs_dat_i[10] wbs_dat_i[11] wbs_dat_i[12] wbs_dat_i[13]
+ wbs_dat_i[14] wbs_dat_i[15] wbs_dat_i[16] wbs_dat_i[17] wbs_dat_i[18] wbs_dat_i[19]
+ wbs_dat_i[1] wbs_dat_i[20] wbs_dat_i[21] wbs_dat_i[22] wbs_dat_i[23] wbs_dat_i[24]
+ wbs_dat_i[25] wbs_dat_i[26] wbs_dat_i[27] wbs_dat_i[28] wbs_dat_i[29] wbs_dat_i[2]
+ wbs_dat_i[30] wbs_dat_i[31] wbs_dat_i[3] wbs_dat_i[4] wbs_dat_i[5] wbs_dat_i[6]
+ wbs_dat_i[7] wbs_dat_i[8] wbs_dat_i[9] wbs_dat_o[0] wbs_dat_o[10] wbs_dat_o[11]
+ wbs_dat_o[12] wbs_dat_o[13] wbs_dat_o[14] wbs_dat_o[15] wbs_dat_o[16] wbs_dat_o[17]
+ wbs_dat_o[18] wbs_dat_o[19] wbs_dat_o[1] wbs_dat_o[20] wbs_dat_o[21] wbs_dat_o[22]
+ wbs_dat_o[23] wbs_dat_o[24] wbs_dat_o[25] wbs_dat_o[26] wbs_dat_o[27] wbs_dat_o[28]
+ wbs_dat_o[29] wbs_dat_o[2] wbs_dat_o[30] wbs_dat_o[31] wbs_dat_o[3] wbs_dat_o[4]
+ wbs_dat_o[5] wbs_dat_o[6] wbs_dat_o[7] wbs_dat_o[8] wbs_dat_o[9] wbs_sel_i[0] wbs_sel_i[1]
+ wbs_sel_i[2] wbs_sel_i[3] wbs_stb_i wbs_we_i
XFILLER_67_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3155_ soc.spi_video_ram_1.buffer_index\[5\] _0769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_82_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3086_ _0705_ _0706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_27_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3988_ _1510_ _1550_ _1551_ _0033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6776_ _0618_ clknet_leaf_84_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[1\]\[18\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5727_ _2817_ _0506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xcaravel_hack_soc_229 io_oeb[33] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
X_5658_ _0878_ _2778_ _2780_ _0474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xcaravel_hack_soc_218 wbs_dat_o[25] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xcaravel_hack_soc_207 wbs_dat_o[14] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_123_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4609_ soc.spi_video_ram_1.write_fifo.fifo_mem\[4\]\[0\] soc.spi_video_ram_1.fifo_in_data\[0\]
+ _2058_ _2059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5589_ soc.spi_video_ram_1.fifo_in_address\[10\] soc.spi_video_ram_1.write_fifo.fifo_mem\[5\]\[26\]
+ _2719_ _2735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_117_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_78_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1800 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1822 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1833 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1811 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1866 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1855 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1844 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1899 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1888 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1877 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_60_wb_clk_i clknet_4_13_0_wb_clk_i clknet_leaf_60_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_77_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4960_ _2290_ _0266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4891_ soc.rom_encoder_0.input_buffer\[2\] _2247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3911_ _1410_ _1439_ _1477_ _1480_ _1484_ _1485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_44_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6630_ soc.cpu.PC.in\[13\] net87 soc.cpu.AReg.data\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_3842_ _1425_ _1428_ _1429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_20_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6561_ _0434_ clknet_leaf_82_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[5\]\[9\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_34_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5512_ _0675_ _2690_ _2691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_3773_ _0760_ _0830_ _1365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6492_ _0365_ clknet_leaf_61_wb_clk_i soc.ram_encoder_0.request_data_out\[5\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_105_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5443_ soc.ram_data_out\[8\] _2603_ _2639_ _2640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_114_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5374_ soc.ram_encoder_0.address\[9\] soc.ram_encoder_0.request_address\[9\] _2581_
+ _2586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_114_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4325_ _1129_ _1851_ _0729_ _1852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_114_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4256_ soc.spi_video_ram_1.write_fifo.fifo_mem\[5\]\[8\] _1787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_83_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3207_ _0757_ soc.spi_video_ram_1.output_buffer\[23\] _0821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4187_ soc.spi_video_ram_1.write_fifo.fifo_mem\[0\]\[3\] soc.spi_video_ram_1.write_fifo.fifo_mem\[1\]\[3\]
+ soc.spi_video_ram_1.write_fifo.fifo_mem\[2\]\[3\] soc.spi_video_ram_1.write_fifo.fifo_mem\[3\]\[3\]
+ _1585_ _1711_ _1723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_95_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3138_ soc.spi_video_ram_1.buffer_index\[3\] _0752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_27_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3069_ net18 _0689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_6828_ _0670_ clknet_leaf_50_wb_clk_i soc.ram_encoder_0.data_out\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_50_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6759_ _0601_ clknet_leaf_126_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[1\]\[1\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_124_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xcaravel_hack_soc_94 io_oeb[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_18_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1696 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_128_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4110_ soc.cpu.AReg.data\[15\] _1658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5090_ _2375_ _0311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_25_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_111_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4041_ _1596_ _1597_ _1598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_65_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5992_ _2985_ _2988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_4943_ _2281_ _0258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_32_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6613_ _0470_ clknet_leaf_20_wb_clk_i soc.rom_loader.current_address\[13\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_71_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4874_ _1426_ _2234_ _2235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3825_ soc.rom_encoder_0.current_state\[2\] _1408_ _1412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_21_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6544_ _0417_ clknet_leaf_41_wb_clk_i soc.ram_encoder_0.initializing_step\[4\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_119_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3756_ _1126_ _1127_ _1167_ _1211_ _1354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_134_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6475_ _0348_ clknet_leaf_58_wb_clk_i soc.ram_encoder_0.input_buffer\[1\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5426_ _2502_ _2624_ _2625_ _2626_ _2627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_3687_ _1278_ _1282_ _1283_ _1284_ _1285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_5357_ soc.ram_encoder_0.address\[1\] soc.ram_encoder_0.request_address\[1\] _2566_
+ _2577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5288_ _2526_ _2505_ _2527_ _0357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_99_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4308_ _1257_ _1835_ _1836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_114_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4239_ _1596_ _1770_ _1771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_28_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_124_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_111_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2150 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2161 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2183 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2172 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4590_ soc.spi_video_ram_1.fifo_in_address\[5\] soc.spi_video_ram_1.write_fifo.fifo_mem\[7\]\[21\]
+ _2037_ _2048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3610_ _1196_ _1197_ _1207_ _1208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_30_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3541_ soc.video_generator_1.v_count\[0\] _1139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_143_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3472_ _0907_ soc.cpu.AReg.data\[12\] _1012_ soc.ram_data_out\[12\] _1073_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6260_ _0135_ clknet_leaf_83_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[7\]\[18\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_142_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5211_ _1413_ _2465_ _2470_ _0337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6191_ _0071_ clknet_leaf_116_wb_clk_i soc.spi_video_ram_1.output_buffer\[9\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_43_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5142_ _2400_ _2417_ _0321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_96_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5073_ _2366_ _0303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_84_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4024_ _1580_ _1581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_93_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5975_ soc.spi_video_ram_1.write_fifo.fifo_mem\[0\]\[23\] soc.spi_video_ram_1.fifo_in_address\[7\]
+ _2952_ _2978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4926_ _2271_ _2272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_52_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4857_ _1461_ _1953_ _1954_ _0234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_119_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3808_ _1379_ _1393_ _1398_ _1386_ _1399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_6527_ _0400_ clknet_leaf_57_wb_clk_i soc.ram_data_out\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4788_ _0720_ _2176_ _2177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3739_ _1167_ _1336_ _1337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6458_ _0331_ clknet_leaf_16_wb_clk_i soc.cpu.instruction\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_133_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5409_ _2604_ _2611_ _2612_ _2613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_6389_ _0262_ clknet_leaf_24_wb_clk_i soc.rom_encoder_0.request_data_out\[10\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_102_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_48_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_117_wb_clk_i clknet_4_8_0_wb_clk_i clknet_leaf_117_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_44_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_129_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_109_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5760_ _0958_ _0970_ _1002_ _2835_ _2836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_15_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4711_ _2118_ _0189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5691_ _2797_ _2798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_4642_ soc.spi_video_ram_1.write_fifo.fifo_mem\[4\]\[16\] soc.spi_video_ram_1.fifo_in_address\[0\]
+ _2069_ _2076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_116_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4573_ _2039_ _0129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_144_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3524_ _0990_ _1122_ _1123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_6312_ _0187_ clknet_leaf_140_wb_clk_i soc.spi_video_ram_1.sram_sck_fall_edge vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_115_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3455_ _0990_ _1057_ _1058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_6243_ _0118_ clknet_leaf_126_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[7\]\[1\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_118_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6174_ _0054_ clknet_leaf_67_wb_clk_i soc.ram_encoder_0.output_buffer\[3\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3386_ _0979_ _0984_ soc.cpu.ALU.f _0986_ _0992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_58_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5125_ soc.cpu.DMuxJMP.sel\[1\] _2392_ _2403_ _2404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_69_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5056_ soc.spi_video_ram_1.write_fifo.fifo_mem\[3\]\[8\] soc.spi_video_ram_1.fifo_in_data\[8\]
+ _2357_ _2358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_38_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4007_ soc.ram_encoder_0.output_buffer\[17\] _1527_ _1568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_66_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_53_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5958_ _2969_ _0585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_41_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4909_ _2258_ _2242_ _2259_ _0246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_21_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5889_ soc.boot_loading_offset\[3\] _2925_ _2927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_138_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_85_wb_clk_i clknet_4_9_0_wb_clk_i clknet_leaf_85_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
Xclkbuf_leaf_14_wb_clk_i clknet_4_3_0_wb_clk_i clknet_leaf_14_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_6_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3240_ soc.cpu.ALU.ny _0853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XTAP_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3171_ soc.spi_video_ram_1.output_buffer\[9\] soc.spi_video_ram_1.output_buffer\[8\]
+ _0783_ _0785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_35_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5812_ soc.cpu.PC.REG.data\[8\] soc.cpu.PC.REG.data\[9\] _2872_ _2878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_63_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6792_ _0634_ clknet_leaf_128_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[2\]\[5\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5743_ _2825_ _0514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_22_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5674_ soc.cpu.ALU.x\[8\] _2784_ _2789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_30_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4625_ soc.spi_video_ram_1.write_fifo.fifo_mem\[4\]\[8\] soc.spi_video_ram_1.fifo_in_data\[8\]
+ _2058_ _2067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4556_ _2030_ _0121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3507_ _0972_ _1101_ _1104_ _1106_ _1107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_143_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4487_ _1984_ _1988_ _1989_ _0093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_3438_ _0904_ soc.cpu.ALU.x\[10\] _1041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6226_ _0101_ clknet_leaf_15_wb_clk_i soc.spi_video_ram_1.fifo_in_data\[0\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_6157_ _0037_ clknet_leaf_59_wb_clk_i soc.ram_encoder_0.output_buffer\[18\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3369_ _0887_ soc.cpu.AReg.data\[6\] _0894_ _0976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5108_ _1434_ _1421_ _2388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_57_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6088_ soc.spi_video_ram_1.write_fifo.fifo_mem\[2\]\[17\] soc.spi_video_ram_1.fifo_in_address\[1\]
+ _3031_ _3039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_58_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5039_ soc.spi_video_ram_1.write_fifo.fifo_mem\[3\]\[0\] soc.spi_video_ram_1.fifo_in_data\[0\]
+ _2217_ _2349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_39_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_139_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xoutput75 net75 io_out[28] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput64 net64 io_out[16] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput53 net53 io_oeb[19] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_110_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_132_wb_clk_i clknet_4_2_0_wb_clk_i clknet_leaf_132_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_88_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4410_ _1585_ _1930_ _1931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_8_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5390_ _1495_ _2595_ _2596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_125_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4341_ _1593_ _1866_ _1867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_114_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4272_ _1711_ _1798_ _1801_ _1761_ _1802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_28_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6011_ soc.spi_video_ram_1.fifo_in_data\[10\] soc.spi_video_ram_1.write_fifo.fifo_mem\[1\]\[10\]
+ _2986_ _2998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3223_ _0776_ soc.spi_video_ram_1.output_buffer\[1\] _0759_ _0837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_39_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3154_ _0767_ _0768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_55_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3085_ soc.spi_video_ram_1.current_state\[3\] soc.spi_video_ram_1.current_state\[0\]
+ _0704_ _0705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_54_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_22_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3987_ soc.ram_encoder_0.output_buffer\[14\] _1527_ _1551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6775_ _0617_ clknet_leaf_74_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[1\]\[17\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5726_ soc.spi_video_ram_1.write_fifo.fifo_mem\[6\]\[16\] soc.spi_video_ram_1.fifo_in_address\[0\]
+ _2810_ _2817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_10_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xcaravel_hack_soc_208 wbs_dat_o[15] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xcaravel_hack_soc_219 wbs_dat_o[26] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_5657_ soc.cpu.ALU.x\[0\] _2779_ _2780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5588_ _2734_ _0450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4608_ _2057_ _2058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_116_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4539_ soc.spi_video_ram_1.fifo_in_data\[14\] _2018_ _2020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6209_ _0084_ clknet_leaf_139_wb_clk_i soc.spi_video_ram_1.state_counter\[4\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_131_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_73_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1823 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1834 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1801 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1867 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1856 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1889 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1878 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_96_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_114_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_64_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4890_ _2245_ _2242_ _2246_ _0240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3910_ soc.rom_encoder_0.request_data_out\[12\] _1481_ _1482_ soc.rom_encoder_0.output_buffer\[16\]
+ _1483_ _1484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_3841_ _1406_ _1427_ _1428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_20_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3772_ _0749_ _1363_ _1364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_34_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6560_ _0433_ clknet_leaf_121_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[5\]\[8\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5511_ _2686_ soc.hack_clock_0.counter\[1\] _2688_ _2689_ _2690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_73_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6491_ _0364_ clknet_leaf_63_wb_clk_i soc.ram_encoder_0.request_data_out\[4\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5442_ _2514_ _2624_ _2625_ _2638_ _2639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_5373_ _2585_ _0384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4324_ _1127_ _1167_ _1851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_87_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4255_ _1596_ _1784_ _1785_ _1786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_110_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3206_ soc.spi_video_ram_1.output_buffer\[22\] _0820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4186_ _1715_ _1686_ _1721_ _1722_ _0059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_41_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3137_ _0750_ soc.spi_video_ram_1.buffer_index\[1\] _0751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_27_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3068_ _0676_ _0688_ _0003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6827_ _0669_ clknet_leaf_48_wb_clk_i soc.ram_encoder_0.data_out\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_50_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6758_ _0600_ clknet_leaf_10_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[1\]\[0\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_6_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6689_ _0531_ net84 soc.cpu.PC.REG.data\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5709_ soc.spi_video_ram_1.write_fifo.fifo_mem\[6\]\[8\] soc.spi_video_ram_1.fifo_in_data\[8\]
+ _2799_ _2808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_136_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xcaravel_hack_soc_95 io_oeb[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_15_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_42_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1697 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_4_12_0_wb_clk_i clknet_0_wb_clk_i clknet_4_12_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_4040_ soc.spi_video_ram_1.write_fifo.fifo_mem\[5\]\[16\] _1597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_64_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5991_ _2987_ _0600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_80_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4942_ soc.rom_encoder_0.data_out\[6\] soc.rom_encoder_0.request_data_out\[6\] _2276_
+ _2281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6612_ _0469_ clknet_leaf_20_wb_clk_i soc.rom_loader.current_address\[12\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4873_ soc.rom_encoder_0.input_bits_left\[2\] _2232_ _2234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_21_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3824_ soc.rom_encoder_0.request_write _1411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_32_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6543_ _0416_ clknet_leaf_34_wb_clk_i soc.ram_encoder_0.initializing_step\[3\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3755_ _1142_ soc.video_generator_1.v_count\[7\] _1353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_6474_ _0347_ clknet_leaf_45_wb_clk_i soc.ram_encoder_0.input_buffer\[0\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3686_ _1272_ _1239_ _1266_ _1284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_118_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5425_ soc.ram_encoder_0.request_data_out\[4\] _2606_ _2626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_142_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_114_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5356_ _2576_ _0376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5287_ soc.ram_encoder_0.input_buffer\[6\] _2503_ _2508_ _2527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_101_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4307_ _1127_ _1167_ _1835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_75_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4238_ soc.spi_video_ram_1.write_fifo.fifo_mem\[7\]\[7\] _1770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_68_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_67_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4169_ _1595_ soc.spi_video_ram_1.write_fifo.fifo_mem\[4\]\[1\] _1706_ _1707_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_71_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_3_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xclkbuf_leaf_39_wb_clk_i clknet_4_7_0_wb_clk_i clknet_leaf_39_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_78_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2151 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2162 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2140 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2184 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2173 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3540_ soc.ram_encoder_0.initialized soc.spi_video_ram_1.initialized _1137_ _1138_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_31_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_142_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3471_ _0923_ _1071_ _1072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_5210_ _1426_ _2468_ _1428_ _0690_ _2470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_130_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6190_ _0070_ clknet_leaf_116_wb_clk_i soc.spi_video_ram_1.output_buffer\[10\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_124_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5141_ soc.cpu.instruction\[4\] _2392_ _2416_ _2417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_36_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5072_ soc.spi_video_ram_1.write_fifo.fifo_mem\[3\]\[16\] soc.spi_video_ram_1.fifo_in_address\[0\]
+ _2357_ _2366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_96_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4023_ _1579_ _1580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_65_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5974_ _2977_ _0593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_100_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4925_ _2270_ _2271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
X_4856_ _1461_ _1951_ _1952_ _0233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_3807_ _1383_ _1394_ _1397_ _1379_ _1398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_6526_ _0399_ clknet_leaf_55_wb_clk_i soc.ram_data_out\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4787_ _0674_ soc.spi_video_ram_1.sram_sck_rise_edge _2176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_134_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3738_ _1162_ soc.video_generator_1.v_count\[2\] _1336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6457_ _0330_ clknet_leaf_19_wb_clk_i soc.cpu.instruction\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3669_ _1218_ _1266_ _1261_ _1267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5408_ net2 _2488_ _2612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6388_ _0261_ clknet_leaf_36_wb_clk_i soc.rom_encoder_0.request_data_out\[9\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5339_ soc.ram_encoder_0.data_out\[11\] _2565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_88_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_12_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_8_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_125_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_120_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4710_ net9 soc.spi_video_ram_1.read_value\[0\] _2117_ _2118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5690_ _0700_ _2703_ _0698_ _2797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_4641_ _2075_ _0161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_30_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_129_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_116_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4572_ soc.spi_video_ram_1.fifo_in_data\[12\] soc.spi_video_ram_1.write_fifo.fifo_mem\[7\]\[12\]
+ _2037_ _2039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_143_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3523_ _0972_ _1116_ _1120_ _1121_ _1122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
X_6311_ _0186_ clknet_leaf_135_wb_clk_i soc.spi_video_ram_1.sram_sck_rise_edge vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_7_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_144_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3454_ _0972_ _1054_ _1055_ _1056_ _1057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_6242_ _0117_ clknet_leaf_12_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[7\]\[0\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_131_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6173_ _0053_ clknet_leaf_65_wb_clk_i soc.ram_encoder_0.output_buffer\[4\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_97_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3385_ _0884_ _0989_ _0991_ soc.cpu.PC.in\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_112_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5124_ _2393_ _2401_ _2402_ _2403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_69_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5055_ _2216_ _2357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_4006_ _1557_ _1559_ _1566_ _1567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_84_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5957_ soc.spi_video_ram_1.write_fifo.fifo_mem\[0\]\[14\] soc.spi_video_ram_1.fifo_in_data\[14\]
+ _2964_ _2969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_139_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4908_ soc.rom_encoder_0.input_buffer\[3\] _2243_ _2250_ _2259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_40_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5888_ soc.boot_loading_offset\[3\] _2925_ _2926_ _0558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_21_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4839_ soc.spi_video_ram_1.initialized soc.video_generator_1.h_count\[1\] _1189_
+ _2207_ _2208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_135_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6509_ _0382_ clknet_leaf_67_wb_clk_i soc.ram_encoder_0.request_address\[6\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_106_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_76_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_91_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_54_wb_clk_i clknet_4_12_0_wb_clk_i clknet_leaf_54_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_141_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3170_ soc.spi_video_ram_1.output_buffer\[11\] soc.spi_video_ram_1.output_buffer\[10\]
+ _0783_ _0784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_66_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_82_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5811_ _2847_ _2876_ _2877_ _2849_ _0529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_62_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6791_ _0633_ clknet_leaf_9_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[2\]\[4\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5742_ soc.spi_video_ram_1.write_fifo.fifo_mem\[6\]\[24\] soc.spi_video_ram_1.fifo_in_address\[8\]
+ _2798_ _2825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5673_ _1002_ _2778_ _2788_ _0481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_30_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4624_ _2066_ _0153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4555_ soc.spi_video_ram_1.fifo_in_data\[4\] soc.spi_video_ram_1.write_fifo.fifo_mem\[7\]\[4\]
+ _2023_ _2030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_144_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3506_ _0972_ _1105_ _1106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4486_ soc.video_generator_1.v_count\[2\] _1987_ _1989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_104_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3437_ _0884_ _1039_ _1040_ soc.cpu.PC.in\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_6225_ _0100_ clknet_leaf_141_wb_clk_i soc.video_generator_1.v_count\[9\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6156_ _0036_ clknet_leaf_60_wb_clk_i soc.ram_encoder_0.output_buffer\[17\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_98_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3368_ soc.ram_data_out\[6\] _0869_ _0868_ net43 _0854_ _0975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_44_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5107_ _0691_ _2387_ _0316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3299_ net79 _0855_ _0860_ _0862_ _0910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
X_6087_ _3038_ _0645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_57_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5038_ _2330_ _2347_ _2348_ _0676_ _0286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_73_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_25_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_53_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xoutput65 net65 io_out[17] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput76 net76 io_out[29] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput54 net54 io_oeb[22] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xclkbuf_leaf_101_wb_clk_i clknet_4_10_0_wb_clk_i clknet_leaf_101_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_44_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_108_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_8_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4340_ soc.spi_video_ram_1.write_fifo.fifo_mem\[5\]\[13\] _1866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_4_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4271_ _1756_ _1799_ _1800_ _1710_ _1801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_140_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6010_ _1799_ _2988_ _2997_ _0609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3222_ _0835_ _0836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_79_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3153_ soc.spi_video_ram_1.output_buffer\[1\] _0763_ _0765_ _0766_ _0767_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_55_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3084_ _0703_ soc.spi_video_ram_1.current_state\[4\] _0704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_39_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3986_ soc.ram_encoder_0.output_buffer\[10\] _1520_ _1530_ soc.ram_encoder_0.request_data_out\[6\]
+ _1549_ _1550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_6774_ _0616_ clknet_leaf_79_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[1\]\[16\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5725_ _2816_ _0505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_22_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5656_ _2777_ _2779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_30_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4607_ _2056_ _2057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
Xcaravel_hack_soc_209 wbs_dat_o[16] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_11_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5587_ soc.spi_video_ram_1.fifo_in_address\[9\] soc.spi_video_ram_1.write_fifo.fifo_mem\[5\]\[25\]
+ _2719_ _2734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_105_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4538_ _2003_ _1108_ _2019_ _0114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_144_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4469_ _1960_ _1975_ _1976_ _0088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_77_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6208_ _0083_ clknet_leaf_139_wb_clk_i soc.spi_video_ram_1.state_counter\[3\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_100_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6139_ _0019_ clknet_leaf_1_wb_clk_i soc.video_generator_1.h_count\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_85_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_46_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1824 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1813 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1802 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1857 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1846 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1835 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1879 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1868 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_36_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3840_ _1426_ soc.rom_encoder_0.current_state\[1\] _1427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_3771_ _0758_ _0759_ _0752_ _1363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_20_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5510_ soc.hack_clock_0.counter\[3\] soc.hack_clock_0.counter\[2\] _2689_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6490_ _0363_ clknet_leaf_63_wb_clk_i soc.ram_encoder_0.request_data_out\[3\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_9_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5441_ soc.ram_encoder_0.request_data_out\[8\] _2605_ _2638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_66_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5372_ soc.ram_encoder_0.address\[8\] soc.ram_encoder_0.request_address\[8\] _2581_
+ _2585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_114_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4323_ _0703_ _0686_ _1850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_141_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4254_ _1600_ soc.spi_video_ram_1.write_fifo.fifo_mem\[2\]\[8\] _1587_ _1785_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_101_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3205_ _0752_ _0818_ _0819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4185_ _0720_ _1692_ _1578_ _1696_ _1722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_83_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3136_ soc.spi_video_ram_1.buffer_index\[0\] _0750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_3067_ soc.spi_video_ram_1.current_state\[0\] _0687_ _0688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_43_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6826_ _0668_ clknet_leaf_48_wb_clk_i soc.ram_encoder_0.data_out\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_50_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6757_ _0599_ clknet_leaf_110_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[0\]\[28\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_23_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3969_ soc.ram_encoder_0.request_address\[9\] _1513_ _1537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_50_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5708_ _2807_ _0497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_137_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6688_ _0530_ net85 soc.cpu.PC.REG.data\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_12_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5639_ _2746_ _2766_ _2767_ _0467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_144_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xcaravel_hack_soc_96 io_oeb[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_2344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1698 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5990_ soc.spi_video_ram_1.fifo_in_data\[0\] soc.spi_video_ram_1.write_fifo.fifo_mem\[1\]\[0\]
+ _2986_ _2987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_25_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4941_ _2280_ _0257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_17_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4872_ soc.rom_encoder_0.input_bits_left\[2\] _2232_ _2233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6611_ _0468_ clknet_leaf_20_wb_clk_i soc.rom_loader.current_address\[11\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3823_ _1406_ _1409_ _1410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_119_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6542_ _0415_ clknet_leaf_34_wb_clk_i soc.ram_encoder_0.initializing_step\[2\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_3754_ _1142_ soc.video_generator_1.v_count\[8\] _1352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xclkbuf_leaf_9_wb_clk_i clknet_4_1_0_wb_clk_i clknet_leaf_9_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_6473_ _0346_ clknet_leaf_41_wb_clk_i soc.ram_encoder_0.input_bits_left\[4\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_119_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3685_ _1272_ _1239_ _1270_ _1283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5424_ _2602_ _2625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_5355_ soc.ram_encoder_0.address\[0\] soc.ram_encoder_0.request_address\[0\] _2566_
+ _2576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_99_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5286_ soc.ram_encoder_0.input_buffer\[10\] _2526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_102_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4306_ _1609_ _1833_ _1834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4237_ _1595_ soc.spi_video_ram_1.write_fifo.fifo_mem\[4\]\[7\] _1768_ _1769_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_96_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_74_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4168_ _1596_ _1705_ _1706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_83_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4099_ _1414_ _1647_ _1649_ _1646_ _0045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_56_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3119_ _0708_ _0702_ _0706_ _0736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_55_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_24_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6809_ _0651_ clknet_leaf_98_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[2\]\[22\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_11_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_93_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_47_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_79_wb_clk_i clknet_4_14_0_wb_clk_i clknet_leaf_79_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_46_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2152 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2141 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2130 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2185 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2174 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2163 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_11_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3470_ _0904_ soc.cpu.ALU.x\[12\] _1071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_7_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_142_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5140_ _2240_ _2413_ _2414_ _2415_ _2416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_97_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5071_ _2365_ _0302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_29_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_56_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4022_ _0002_ _1579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_38_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5973_ soc.spi_video_ram_1.write_fifo.fifo_mem\[0\]\[22\] soc.spi_video_ram_1.fifo_in_address\[6\]
+ _2952_ _2977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4924_ _1403_ _0674_ _2268_ _2269_ _2270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_21_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4855_ _0691_ _2219_ _0232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4786_ _1671_ _2174_ _2175_ _0207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3806_ _1383_ _1395_ _1396_ _1397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_20_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6525_ _0398_ clknet_leaf_58_wb_clk_i soc.ram_data_out\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3737_ _1333_ _1242_ _1208_ _1334_ _1335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_118_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_106_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6456_ _0329_ clknet_leaf_48_wb_clk_i soc.cpu.instruction\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3668_ soc.video_generator_1.h_count\[2\] _1217_ _1266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_134_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5407_ soc.ram_encoder_0.request_data_out\[1\] _2606_ _2611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6387_ _0260_ clknet_leaf_11_wb_clk_i soc.rom_encoder_0.request_data_out\[8\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3599_ soc.video_generator_1.h_count\[3\] soc.video_generator_1.h_count\[4\] _1196_
+ _1197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_5338_ _2563_ _2538_ _2564_ _0370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_134_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_130_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5269_ soc.ram_encoder_0.input_buffer\[0\] _2505_ _2508_ _2515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_75_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xclkbuf_leaf_126_wb_clk_i clknet_4_3_0_wb_clk_i clknet_leaf_126_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_137_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4640_ soc.spi_video_ram_1.write_fifo.fifo_mem\[4\]\[15\] soc.spi_video_ram_1.fifo_in_data\[15\]
+ _2069_ _2075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_144_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4571_ _2038_ _0128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6310_ _0185_ clknet_leaf_138_wb_clk_i net69 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
X_3522_ _0972_ _1111_ _1114_ _1121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_7_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3453_ _0972_ _1042_ _1045_ _1056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_6241_ _0116_ clknet_leaf_75_wb_clk_i soc.spi_video_ram_1.fifo_in_data\[15\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_143_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6172_ _0052_ clknet_leaf_26_wb_clk_i soc.rom_encoder_0.output_buffer\[1\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3384_ _0846_ _0990_ soc.cpu.AReg.data\[6\] _0881_ _0991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_5123_ net6 _2223_ _2402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_58_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5054_ _2356_ _0294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4005_ _1563_ _1565_ _1566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_84_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5956_ _2968_ _0584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_34_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4907_ soc.rom_encoder_0.input_buffer\[7\] _2258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5887_ soc.boot_loading_offset\[3\] _2925_ _0675_ _2926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4838_ _1216_ _1131_ _2206_ _2207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_14_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4769_ soc.rom_encoder_0.output_buffer\[16\] _2138_ _2162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_5_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6508_ _0381_ clknet_leaf_66_wb_clk_i soc.ram_encoder_0.request_address\[5\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_20_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_135_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6439_ _0312_ clknet_leaf_109_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[3\]\[25\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_106_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_32_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_94_wb_clk_i clknet_4_11_0_wb_clk_i clknet_leaf_94_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xclkbuf_leaf_23_wb_clk_i clknet_4_4_0_wb_clk_i clknet_leaf_23_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_39_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5810_ soc.cpu.PC.in\[9\] _2851_ _2877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_35_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6790_ _0632_ clknet_leaf_9_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[2\]\[3\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_96_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5741_ _2824_ _0513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_16_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5672_ soc.cpu.ALU.x\[7\] _2784_ _2788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_135_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4623_ soc.spi_video_ram_1.write_fifo.fifo_mem\[4\]\[7\] soc.spi_video_ram_1.fifo_in_data\[7\]
+ _2058_ _2066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_129_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4554_ _2029_ _0120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_144_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3505_ _1096_ _1099_ _1105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_144_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6224_ _0099_ clknet_leaf_140_wb_clk_i soc.video_generator_1.v_count\[8\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_4485_ soc.video_generator_1.v_count\[2\] _1987_ _1988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_131_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3436_ _0845_ _1011_ soc.cpu.AReg.data\[9\] _0880_ _1040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_6155_ _0035_ clknet_leaf_44_wb_clk_i soc.ram_encoder_0.output_buffer\[16\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_106_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3367_ _0849_ _0973_ _0974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6086_ soc.spi_video_ram_1.write_fifo.fifo_mem\[2\]\[16\] soc.spi_video_ram_1.fifo_in_address\[0\]
+ _3031_ _3038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5106_ soc.rom_encoder_0.initialized _2386_ _2387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5037_ net61 _2330_ _2348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3298_ soc.ram_data_out\[2\] _0869_ _0854_ _0909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_85_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_25_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_41_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5939_ _2959_ _0576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_21_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput55 net55 io_oeb[23] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput66 net66 io_out[18] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_1_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xoutput77 net77 io_out[34] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_141_wb_clk_i clknet_4_2_0_wb_clk_i clknet_leaf_141_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XPHY_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_8_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_117_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_67_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4270_ _1724_ soc.spi_video_ram_1.write_fifo.fifo_mem\[0\]\[9\] _1800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_97_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3221_ _0757_ _0833_ _0834_ _0759_ _0835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_100_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3152_ soc.spi_video_ram_1.output_buffer\[3\] soc.spi_video_ram_1.output_buffer\[2\]
+ _0750_ _0766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_95_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_67_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3083_ soc.spi_video_ram_1.current_state\[1\] _0703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_27_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3985_ soc.ram_encoder_0.request_address\[13\] _1513_ _1549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_6773_ _0615_ clknet_leaf_72_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[1\]\[15\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_50_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5724_ soc.spi_video_ram_1.write_fifo.fifo_mem\[6\]\[15\] soc.spi_video_ram_1.fifo_in_data\[15\]
+ _2810_ _2816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_109_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5655_ _2777_ _2778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_4606_ _0700_ _0694_ _0698_ _2056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_5586_ _2733_ _0449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_144_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4537_ soc.spi_video_ram_1.fifo_in_data\[13\] _2018_ _2019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_117_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4468_ soc.spi_video_ram_1.state_counter\[8\] _1973_ _1976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3419_ _0922_ _1023_ _1024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_6207_ _0082_ clknet_leaf_139_wb_clk_i soc.spi_video_ram_1.state_counter\[2\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_86_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_58_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4399_ _1695_ _1921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6138_ _0018_ clknet_leaf_1_wb_clk_i soc.video_generator_1.h_count\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6069_ soc.spi_video_ram_1.write_fifo.fifo_mem\[2\]\[8\] soc.spi_video_ram_1.fifo_in_data\[8\]
+ _3020_ _3029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_54_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1825 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1814 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1803 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1858 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1847 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1836 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1869 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_10_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_123_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_91_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_44_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_33_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3770_ _0752_ _0808_ _1362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_118_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5440_ _2615_ _2637_ _0399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_9_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5371_ _2584_ _0383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_59_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4322_ _1702_ _1845_ _1848_ _1849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_114_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4253_ soc.spi_video_ram_1.write_fifo.fifo_mem\[3\]\[8\] _1784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_101_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3204_ _0813_ _0817_ _0818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4184_ _1581_ _1716_ _1719_ _1720_ _1721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_68_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3135_ soc.spi_video_ram_1.buffer_index\[4\] _0749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_94_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3066_ _0680_ _0686_ _0687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_70_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6825_ _0667_ clknet_leaf_48_wb_clk_i soc.ram_encoder_0.data_out\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_24_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3968_ _1510_ _1535_ _1536_ _0028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_23_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6756_ _0598_ clknet_leaf_101_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[0\]\[27\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5707_ soc.spi_video_ram_1.write_fifo.fifo_mem\[6\]\[7\] soc.spi_video_ram_1.fifo_in_data\[7\]
+ _2799_ _2807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_136_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6687_ _0529_ net85 soc.cpu.PC.REG.data\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3899_ _1130_ _1472_ _1474_ _0021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5638_ soc.rom_loader.current_address\[10\] _2765_ _2767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_105_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5569_ soc.spi_video_ram_1.fifo_in_address\[0\] _2708_ _2725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_132_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xcaravel_hack_soc_97 io_oeb[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_2334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_139_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_128_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4940_ soc.rom_encoder_0.data_out\[5\] soc.rom_encoder_0.request_data_out\[5\] _2276_
+ _2280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_64_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4871_ _2222_ _2223_ _2231_ _2232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_21_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6610_ _0467_ clknet_leaf_29_wb_clk_i soc.rom_loader.current_address\[10\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3822_ _1407_ _1408_ _1409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_33_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6541_ _0414_ clknet_leaf_34_wb_clk_i soc.ram_encoder_0.initializing_step\[1\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_20_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3753_ _1349_ _1217_ _1218_ _1350_ _1351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_6472_ _0345_ clknet_leaf_41_wb_clk_i soc.ram_encoder_0.input_bits_left\[3\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3684_ _1279_ _1280_ _1281_ _1282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_134_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5423_ _2605_ _2624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_5354_ _2574_ _2538_ _2575_ _0375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_114_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4305_ _1831_ _1832_ _1579_ _1833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_141_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5285_ _2524_ _2504_ _2525_ _0356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_99_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_101_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4236_ _1601_ _1767_ _1768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_114_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_68_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4167_ soc.spi_video_ram_1.write_fifo.fifo_mem\[5\]\[1\] _1705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_95_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3118_ _0703_ _0714_ _0735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4098_ soc.rom_encoder_0.output_bits_left\[2\] _1414_ soc.rom_encoder_0.output_bits_left\[3\]
+ _1648_ _1649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_24_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_142_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6808_ _0650_ clknet_leaf_98_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[2\]\[21\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_51_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6739_ _0581_ clknet_leaf_91_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[0\]\[10\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_20_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_137_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_3_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_2_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2153 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2142 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2131 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2120 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2186 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2175 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2164 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_48_wb_clk_i clknet_4_6_0_wb_clk_i clknet_leaf_48_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_1474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xfanout90 net91 net90 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_70_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_123_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5070_ soc.spi_video_ram_1.write_fifo.fifo_mem\[3\]\[15\] soc.spi_video_ram_1.fifo_in_data\[15\]
+ _2357_ _2365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_111_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4021_ _1577_ _1578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_38_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_80_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5972_ _2976_ _0592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_25_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4923_ soc.hack_rom_request soc.rom_loader.rom_request soc.rom_encoder_0.write_enable
+ _2269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_60_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4854_ _2212_ _2217_ _2218_ _2219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_119_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4785_ soc.rom_encoder_0.output_buffer\[19\] _1670_ _2175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3805_ _0775_ _0773_ _1396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_20_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6524_ _0397_ clknet_leaf_56_wb_clk_i soc.ram_data_out\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3736_ _1142_ soc.video_generator_1.v_count\[7\] _1249_ _1188_ _1334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_106_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6455_ _0328_ clknet_leaf_16_wb_clk_i soc.cpu.ALU.zx vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3667_ _1215_ _1220_ _1265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_115_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5406_ _2436_ _2610_ _0392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6386_ _0259_ clknet_leaf_37_wb_clk_i soc.rom_encoder_0.request_data_out\[7\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3598_ _1133_ _1189_ _1196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_5337_ soc.ram_encoder_0.request_data_out\[10\] _2545_ _2564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_87_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5268_ soc.ram_encoder_0.input_buffer\[4\] _2514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_114_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4219_ _1588_ _1751_ _1752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5199_ _1426_ _1422_ _2459_ _2461_ _0334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_18_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_50_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_79_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_62_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4570_ soc.spi_video_ram_1.fifo_in_data\[11\] soc.spi_video_ram_1.write_fifo.fifo_mem\[7\]\[11\]
+ _2037_ _2038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_30_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3521_ _1117_ _1118_ _1119_ _1120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_144_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3452_ _1049_ _1053_ _1047_ _1055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_6240_ _0115_ clknet_leaf_78_wb_clk_i soc.spi_video_ram_1.fifo_in_data\[14\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_6171_ _0051_ clknet_leaf_26_wb_clk_i soc.rom_encoder_0.output_buffer\[2\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3383_ _0922_ _0990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_69_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xcaravel_hack_soc_190 la_data_out[62] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_41_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5122_ soc.rom_encoder_0.request_data_out\[1\] _2395_ _2401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5053_ soc.spi_video_ram_1.write_fifo.fifo_mem\[3\]\[7\] soc.spi_video_ram_1.fifo_in_data\[7\]
+ _2217_ _2356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_38_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4004_ soc.ram_encoder_0.output_buffer\[13\] _1564_ _1565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_81_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5955_ soc.spi_video_ram_1.write_fifo.fifo_mem\[0\]\[13\] soc.spi_video_ram_1.fifo_in_data\[13\]
+ _2964_ _2968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_80_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4906_ _2256_ _2242_ _2257_ _0245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_40_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5886_ _1461_ _2924_ _2925_ _0557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_4837_ soc.video_generator_1.h_count\[4\] _1132_ _2206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4768_ _1441_ _2160_ _2161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6507_ _0380_ clknet_leaf_65_wb_clk_i soc.ram_encoder_0.request_address\[4\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4699_ soc.spi_video_ram_1.current_state\[2\] net68 _2111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_3719_ _1238_ _1295_ _1316_ _1317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_134_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6438_ _0311_ clknet_leaf_108_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[3\]\[24\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6369_ _0242_ clknet_leaf_19_wb_clk_i soc.rom_encoder_0.input_buffer\[3\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_130_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_76_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_63_wb_clk_i clknet_4_13_0_wb_clk_i clknet_leaf_63_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_63_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5740_ soc.spi_video_ram_1.write_fifo.fifo_mem\[6\]\[23\] soc.spi_video_ram_1.fifo_in_address\[7\]
+ _2798_ _2824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_15_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_89_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5671_ _0989_ _2778_ _2787_ _0480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4622_ _2065_ _0152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_128_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4553_ soc.spi_video_ram_1.fifo_in_data\[3\] soc.spi_video_ram_1.write_fifo.fifo_mem\[7\]\[3\]
+ _2023_ _2029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3504_ _1076_ _1102_ _1103_ _1104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4484_ _1984_ _1986_ _1987_ _0092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_3435_ _0990_ _1038_ _1039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_6223_ _0098_ clknet_leaf_142_wb_clk_i soc.video_generator_1.v_count\[7\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_143_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6154_ _0034_ clknet_leaf_60_wb_clk_i soc.ram_encoder_0.output_buffer\[15\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_98_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3366_ _0850_ soc.cpu.ALU.x\[6\] _0973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3297_ soc.cpu.AReg.data\[2\] _0908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6085_ _3037_ _0644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_58_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5105_ _1438_ _2380_ _2382_ _2385_ _2386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XTAP_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5036_ soc.ram_encoder_0.output_buffer\[19\] _1555_ _1529_ soc.ram_encoder_0.request_data_out\[15\]
+ _1559_ _2347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_100_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_122_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_26_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_54_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5938_ soc.spi_video_ram_1.write_fifo.fifo_mem\[0\]\[5\] soc.spi_video_ram_1.fifo_in_data\[5\]
+ _2953_ _2959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5869_ _2916_ _0549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_22_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput67 net67 io_out[19] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_1_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xoutput56 net56 io_oeb[24] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_89_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput78 net78 io_out[35] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_1_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_131_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_49_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_31_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_leaf_110_wb_clk_i clknet_4_8_0_wb_clk_i clknet_leaf_110_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_114_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_125_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xclkbuf_4_9_0_wb_clk_i clknet_0_wb_clk_i clknet_4_9_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_122_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3220_ _0783_ soc.spi_video_ram_1.output_buffer\[5\] _0834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_79_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3151_ _0751_ _0764_ _0765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_39_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3082_ _0696_ _0699_ _0701_ _0702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_82_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3984_ _1510_ _1547_ _1548_ _0032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_51_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6772_ _0614_ clknet_leaf_88_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[1\]\[14\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_50_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5723_ _2815_ _0504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5654_ _0846_ soc.cpu.instruction\[4\] _2777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_129_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4605_ _2055_ _0145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5585_ soc.spi_video_ram_1.fifo_in_address\[8\] soc.spi_video_ram_1.write_fifo.fifo_mem\[5\]\[24\]
+ _2719_ _2733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_144_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4536_ _0748_ _2018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_131_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4467_ soc.spi_video_ram_1.state_counter\[8\] _1973_ _1975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_3418_ _0875_ _1017_ _1021_ _1022_ _1023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_6206_ _0081_ clknet_leaf_140_wb_clk_i soc.spi_video_ram_1.state_counter\[1\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4398_ _1686_ _1919_ _1920_ _0073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_113_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3349_ _0922_ _0957_ _0958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6137_ _0017_ clknet_leaf_1_wb_clk_i soc.video_generator_1.h_count\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XTAP_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6068_ _3028_ _0636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_39_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5019_ net58 _2330_ _2332_ _2333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_54_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1815 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1804 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_26_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1826 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1837 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_26_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1859 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_111_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5370_ soc.ram_encoder_0.address\[7\] soc.ram_encoder_0.request_address\[7\] _2581_
+ _2584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_113_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4321_ _1580_ _1847_ _1848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_99_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4252_ _1594_ _1781_ _1782_ _1710_ _1783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_3203_ _0760_ _0814_ _0815_ _0816_ _0817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_95_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4183_ _0710_ _1607_ _1720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_41_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3134_ _0748_ _0009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_67_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3065_ _0681_ _0685_ _0686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_82_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6824_ _0666_ clknet_leaf_48_wb_clk_i soc.ram_encoder_0.data_out\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_51_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3967_ soc.ram_encoder_0.output_buffer\[9\] _1527_ _1536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6755_ _0597_ clknet_leaf_103_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[0\]\[26\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5706_ _2806_ _0496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_50_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6686_ _0528_ net85 soc.cpu.PC.REG.data\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3898_ _1462_ _1473_ _1474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5637_ soc.rom_loader.current_address\[10\] _2765_ _2766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_105_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5568_ _2724_ _0440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_105_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4519_ _0009_ _0958_ _2009_ _0105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5499_ soc.ram_encoder_0.initializing_step\[3\] soc.ram_encoder_0.initializing_step\[2\]
+ _2678_ _2680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_132_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_37_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xcaravel_hack_soc_98 io_oeb[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_2335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_77_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_49_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4870_ net18 _2230_ _2231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3821_ soc.rom_encoder_0.current_state\[1\] _1408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_32_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6540_ _0413_ clknet_leaf_35_wb_clk_i soc.ram_encoder_0.initializing_step\[0\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_119_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3752_ soc.spi_video_ram_1.read_value\[0\] _1217_ _1350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6471_ _0344_ clknet_leaf_41_wb_clk_i soc.ram_encoder_0.input_bits_left\[2\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3683_ soc.video_generator_1.h_count\[1\] _1216_ _1281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_5422_ _2615_ _2623_ _0395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5353_ soc.ram_encoder_0.request_data_out\[15\] _2566_ _2575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_126_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4304_ soc.spi_video_ram_1.write_fifo.fifo_mem\[4\]\[27\] soc.spi_video_ram_1.write_fifo.fifo_mem\[5\]\[27\]
+ soc.spi_video_ram_1.write_fifo.fifo_mem\[6\]\[27\] soc.spi_video_ram_1.write_fifo.fifo_mem\[7\]\[27\]
+ _1583_ _1586_ _1832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_5284_ soc.ram_encoder_0.input_buffer\[5\] _2503_ _2508_ _2525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_101_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4235_ soc.spi_video_ram_1.write_fifo.fifo_mem\[5\]\[7\] _1767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4166_ _1700_ _1703_ _1704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_110_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3117_ _0733_ _0734_ _0691_ _0007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4097_ _1478_ _1421_ _1648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_56_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6807_ _0649_ clknet_leaf_119_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[2\]\[20\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4999_ soc.cpu.PC.REG.data\[10\] _2318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_11_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6738_ _0580_ clknet_leaf_122_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[0\]\[9\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_136_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6669_ _0511_ clknet_leaf_97_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[6\]\[21\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_87_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_124_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_19_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2110 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2143 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2132 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2121 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2176 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2154 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2165 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2187 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_42_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_128_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout91 soc.cpu.AReg.clk net91 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_70_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_88_wb_clk_i clknet_4_9_0_wb_clk_i clknet_leaf_88_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_116_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_17_wb_clk_i clknet_4_3_0_wb_clk_i clknet_leaf_17_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_143_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_97_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4020_ _1576_ _0188_ _1577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_37_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_37_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5971_ soc.spi_video_ram_1.write_fifo.fifo_mem\[0\]\[21\] soc.spi_video_ram_1.fifo_in_address\[5\]
+ _2952_ _2976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4922_ soc.rom_encoder_0.current_state\[2\] _1422_ _2268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_127_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4853_ _0694_ _2213_ _0700_ _2218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4784_ soc.rom_encoder_0.output_buffer\[15\] _1436_ _2173_ _1441_ _2174_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_3804_ _0765_ _0777_ _1395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6523_ _0396_ clknet_leaf_56_wb_clk_i soc.ram_data_out\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3735_ _1126_ _1333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_134_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6454_ _0327_ clknet_leaf_51_wb_clk_i soc.cpu.ALU.nx vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_109_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_106_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5405_ soc.ram_data_out\[0\] _2603_ _2609_ _2610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3666_ _1239_ _1263_ _1264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_133_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6385_ _0258_ clknet_leaf_11_wb_clk_i soc.rom_encoder_0.request_data_out\[6\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3597_ _1135_ _1194_ _1195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_130_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5336_ soc.ram_encoder_0.data_out\[10\] _2563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_88_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5267_ _2512_ _2504_ _2513_ _0350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_88_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4218_ soc.spi_video_ram_1.write_fifo.fifo_mem\[0\]\[6\] soc.spi_video_ram_1.write_fifo.fifo_mem\[1\]\[6\]
+ _1724_ _1751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_29_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5198_ soc.rom_encoder_0.sram_sio_oe _2460_ _0690_ _2461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_29_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4149_ soc.spi_video_ram_1.write_fifo.fifo_mem\[4\]\[0\] soc.spi_video_ram_1.write_fifo.fifo_mem\[5\]\[0\]
+ soc.spi_video_ram_1.write_fifo.fifo_mem\[6\]\[0\] soc.spi_video_ram_1.write_fifo.fifo_mem\[7\]\[0\]
+ _1593_ _1587_ _1688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_83_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_54_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_4_11_0_wb_clk_i clknet_0_wb_clk_i clknet_4_11_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_137_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_78_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_135_wb_clk_i clknet_4_2_0_wb_clk_i clknet_leaf_135_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_19_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_91_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_129_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3520_ _1115_ _1119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_144_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_6_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3451_ _1047_ _1049_ _1053_ _1054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_6170_ _0050_ clknet_leaf_26_wb_clk_i soc.rom_encoder_0.output_buffer\[3\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3382_ _0922_ _0988_ _0989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
Xcaravel_hack_soc_191 la_data_out[63] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xcaravel_hack_soc_180 la_data_out[52] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_112_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5121_ _0690_ _2400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_34_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_112_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5052_ _1748_ _2217_ _2355_ _0293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4003_ _1499_ _1515_ _1564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_65_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_80_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_65_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5954_ _2967_ _0583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4905_ soc.rom_encoder_0.input_buffer\[2\] _2243_ _2250_ _2257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_52_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_21_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5885_ soc.boot_loading_offset\[2\] soc.boot_loading_offset\[1\] _2921_ _2925_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_4836_ _2205_ _0227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_21_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6506_ _0379_ clknet_leaf_65_wb_clk_i soc.ram_encoder_0.request_address\[3\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4767_ soc.rom_encoder_0.request_write _1656_ _2158_ _2159_ _2160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_14_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4698_ soc.spi_video_ram_1.state_sram_clk_counter\[7\] _2108_ _2110_ _0183_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3718_ _1310_ _1238_ _1315_ _1316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_6437_ _0310_ clknet_leaf_107_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[3\]\[23\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3649_ _1176_ _1186_ _1246_ _1247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_6368_ _0241_ clknet_leaf_18_wb_clk_i soc.rom_encoder_0.input_buffer\[2\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5319_ soc.ram_encoder_0.request_data_out\[4\] _2545_ _2552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_102_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6299_ _0174_ clknet_leaf_108_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[4\]\[28\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_69_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_57_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xclkbuf_leaf_32_wb_clk_i clknet_4_5_0_wb_clk_i clknet_leaf_32_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_5670_ soc.cpu.ALU.x\[6\] _2784_ _2787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4621_ soc.spi_video_ram_1.write_fifo.fifo_mem\[4\]\[6\] soc.spi_video_ram_1.fifo_in_data\[6\]
+ _2058_ _2065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_117_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4552_ _2028_ _0119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_144_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3503_ _1100_ _1103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_7_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4483_ soc.video_generator_1.v_count\[1\] _1980_ _1987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_3434_ _0972_ _1035_ _1036_ _1037_ _1038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_6222_ _0097_ clknet_leaf_140_wb_clk_i soc.video_generator_1.v_count\[6\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6153_ _0033_ clknet_leaf_62_wb_clk_i soc.ram_encoder_0.output_buffer\[14\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3365_ _0875_ _0972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3296_ _0854_ _0907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_6084_ soc.spi_video_ram_1.write_fifo.fifo_mem\[2\]\[15\] soc.spi_video_ram_1.fifo_in_data\[15\]
+ _3031_ _3037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5104_ soc.rom_encoder_0.initializing_step\[3\] _2383_ _2384_ _2385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5035_ _2330_ _2345_ _2346_ _0676_ _0285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_85_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5937_ _2958_ _0575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_40_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5868_ soc.ram_encoder_0.address\[12\] soc.cpu.AReg.data\[12\] _2902_ _2916_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5799_ _2846_ _2867_ _2868_ _0526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4819_ soc.spi_video_ram_1.fifo_in_address\[4\] soc.cpu.AReg.data\[4\] _2018_ _2197_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_110_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput46 net46 io_oeb[10] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_89_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput57 net57 io_oeb[25] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput79 net79 io_out[36] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_103_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput68 net68 io_out[20] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_130_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_56_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3150_ _0750_ soc.spi_video_ram_1.buffer_index\[1\] _0764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_95_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3081_ soc.spi_video_ram_1.write_fifo.read_pointer\[2\] _0700_ _0701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_36_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6771_ _0613_ clknet_leaf_88_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[1\]\[13\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3983_ soc.ram_encoder_0.output_buffer\[13\] _1527_ _1548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5722_ soc.spi_video_ram_1.write_fifo.fifo_mem\[6\]\[14\] soc.spi_video_ram_1.fifo_in_data\[14\]
+ _2810_ _2815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5653_ soc.rom_loader.wait_fall_clk _2775_ _2776_ _0472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5584_ _2732_ _0448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4604_ soc.spi_video_ram_1.fifo_in_address\[12\] soc.spi_video_ram_1.write_fifo.fifo_mem\[7\]\[28\]
+ _2022_ _2055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4535_ _2003_ _1092_ _2017_ _0113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_7_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4466_ _1961_ _1973_ _1974_ _0087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_3417_ _0875_ _1010_ _1015_ _1022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_6205_ _0080_ clknet_leaf_140_wb_clk_i soc.spi_video_ram_1.state_counter\[0\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4397_ soc.spi_video_ram_1.output_buffer\[7\] _1611_ _1920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_131_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3348_ _0875_ _0953_ _0956_ _0957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6136_ _0016_ clknet_leaf_2_wb_clk_i soc.video_generator_1.h_count\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3279_ net78 _0855_ _0860_ _0862_ _0891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_86_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6067_ soc.spi_video_ram_1.write_fifo.fifo_mem\[2\]\[7\] soc.spi_video_ram_1.fifo_in_data\[7\]
+ _3020_ _3028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_45_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5018_ _2331_ _1508_ _2332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_54_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1816 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1849 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1838 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1827 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_135_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_9_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4320_ _1846_ _1847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_114_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4251_ _1600_ soc.spi_video_ram_1.write_fifo.fifo_mem\[0\]\[8\] _1782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_113_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3202_ soc.spi_video_ram_1.output_buffer\[12\] soc.spi_video_ram_1.output_buffer\[13\]
+ _0783_ _0816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_110_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4182_ _1605_ _1718_ _1719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3133_ _0747_ _0748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_68_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3064_ soc.spi_video_ram_1.state_sram_clk_counter\[8\] soc.spi_video_ram_1.state_sram_clk_counter\[0\]
+ _0684_ _0685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_2
XFILLER_48_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6823_ _0665_ clknet_leaf_56_wb_clk_i soc.ram_encoder_0.data_out\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_50_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_23_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3966_ soc.ram_encoder_0.output_buffer\[5\] _1520_ _1530_ soc.ram_encoder_0.request_data_out\[1\]
+ _1534_ _1535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_6754_ _0596_ clknet_leaf_107_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[0\]\[25\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6685_ _0527_ net84 soc.cpu.PC.REG.data\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5705_ soc.spi_video_ram_1.write_fifo.fifo_mem\[6\]\[6\] soc.spi_video_ram_1.fifo_in_data\[6\]
+ _2799_ _2806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_10_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5636_ _2746_ _2764_ _2765_ _0466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_3897_ _1132_ soc.video_generator_1.h_count\[8\] _1470_ _1473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_128_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5567_ soc.spi_video_ram_1.fifo_in_data\[15\] soc.spi_video_ram_1.write_fifo.fifo_mem\[5\]\[15\]
+ _2719_ _2724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_144_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5498_ soc.ram_encoder_0.initializing_step\[2\] _2678_ _2679_ _0415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4518_ soc.spi_video_ram_1.fifo_in_data\[4\] _2007_ _2009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_2_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4449_ soc.spi_video_ram_1.state_counter\[1\] soc.spi_video_ram_1.state_counter\[0\]
+ soc.spi_video_ram_1.state_counter\[2\] _1963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_144_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6119_ _0970_ _2897_ _3052_ _2553_ _0663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_85_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xcaravel_hack_soc_99 io_oeb[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_27_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_33_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3820_ soc.rom_encoder_0.current_state\[2\] _1407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_3
X_3751_ soc.spi_video_ram_1.read_value\[1\] _1349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6470_ _0343_ clknet_leaf_35_wb_clk_i soc.ram_encoder_0.toggled_sram_sck vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_3682_ _1239_ _1280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_5421_ soc.ram_data_out\[3\] _2603_ _2622_ _2623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_64_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5352_ soc.ram_encoder_0.data_out\[15\] _2574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_114_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4303_ soc.spi_video_ram_1.write_fifo.fifo_mem\[0\]\[27\] soc.spi_video_ram_1.write_fifo.fifo_mem\[1\]\[27\]
+ soc.spi_video_ram_1.write_fifo.fifo_mem\[2\]\[27\] soc.spi_video_ram_1.write_fifo.fifo_mem\[3\]\[27\]
+ _1583_ _1586_ _1831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_142_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5283_ soc.ram_encoder_0.input_buffer\[9\] _2524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_87_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4234_ _0799_ _1686_ _1764_ _1766_ _0063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_67_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4165_ _1592_ _1701_ _1702_ _1703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_110_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3116_ soc.spi_video_ram_1.initialized soc.spi_video_ram_1.start_read soc.spi_video_ram_1.current_state\[2\]
+ _0702_ _0734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_71_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4096_ _1415_ _1646_ _1647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_51_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6806_ _0648_ clknet_leaf_88_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[2\]\[19\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_142_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4998_ _2317_ _0277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_11_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3949_ _1509_ _1522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_6737_ _0579_ clknet_leaf_120_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[0\]\[8\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6668_ _0510_ clknet_leaf_119_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[6\]\[20\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5619_ soc.rom_loader.current_address\[4\] _2753_ _2754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6599_ _0456_ clknet_leaf_7_wb_clk_i soc.rom_encoder_0.toggled_sram_sck vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_136_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_3_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2100 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_73_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2144 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2133 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2122 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2111 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2177 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2155 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2166 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_11_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_6_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_57_wb_clk_i clknet_4_6_0_wb_clk_i clknet_leaf_57_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_97_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_92_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5970_ _2975_ _0591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4921_ _2266_ _2243_ _2267_ _0250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_52_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4852_ _2216_ _2217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_3803_ _0794_ _0796_ _0765_ _1394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4783_ _1413_ _2172_ _2173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6522_ _0395_ clknet_leaf_57_wb_clk_i soc.ram_data_out\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3734_ _1331_ _1150_ _1181_ _1332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_109_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6453_ _0326_ clknet_leaf_51_wb_clk_i soc.cpu.ALU.zy vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3665_ _1241_ _1261_ _1262_ _1263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_118_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5404_ _2604_ _2607_ _2608_ _2609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_115_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6384_ _0257_ clknet_leaf_32_wb_clk_i soc.rom_encoder_0.request_data_out\[5\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_47_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_3596_ soc.video_generator_1.h_count\[5\] _1131_ _1194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_115_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5335_ _2561_ _2538_ _2562_ _0369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_114_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5266_ net4 _2505_ _2508_ _2513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_130_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4217_ _1601_ soc.spi_video_ram_1.write_fifo.fifo_mem\[2\]\[6\] _1749_ _1750_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5197_ _1426_ _2221_ _1424_ _2459_ _2460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or4_1
X_4148_ soc.spi_video_ram_1.write_fifo.fifo_mem\[0\]\[0\] soc.spi_video_ram_1.write_fifo.fifo_mem\[1\]\[0\]
+ soc.spi_video_ram_1.write_fifo.fifo_mem\[2\]\[0\] soc.spi_video_ram_1.write_fifo.fifo_mem\[3\]\[0\]
+ _1594_ _1588_ _1687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_28_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4079_ _1578_ _1632_ _1633_ _0041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_37_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_19_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_104_wb_clk_i clknet_4_10_0_wb_clk_i clknet_leaf_104_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_131_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3450_ _1052_ _1053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_130_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xcaravel_hack_soc_181 la_data_out[53] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_3381_ _0972_ _0985_ _0987_ _0988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xcaravel_hack_soc_192 wbs_ack_o vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xcaravel_hack_soc_170 la_data_out[42] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_5120_ _0691_ _2399_ _0317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5051_ soc.spi_video_ram_1.fifo_in_data\[6\] _2217_ _2355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_27_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4002_ soc.ram_encoder_0.request_data_out\[9\] _1515_ _1529_ _1563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_112_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_38_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_92_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_19_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5953_ soc.spi_video_ram_1.write_fifo.fifo_mem\[0\]\[12\] soc.spi_video_ram_1.fifo_in_data\[12\]
+ _2964_ _2967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_34_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4904_ soc.rom_encoder_0.input_buffer\[6\] _2256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5884_ soc.boot_loading_offset\[1\] _2921_ soc.boot_loading_offset\[2\] _2924_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_139_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4835_ soc.spi_video_ram_1.fifo_in_address\[12\] soc.cpu.AReg.data\[12\] _0748_ _2205_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4766_ soc.rom_encoder_0.request_data_out\[8\] _1481_ _2159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_21_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6505_ _0378_ clknet_leaf_64_wb_clk_i soc.ram_encoder_0.request_address\[2\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3717_ _1280_ _1309_ _1311_ _1314_ _1315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_119_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4697_ soc.spi_video_ram_1.state_sram_clk_counter\[7\] _2108_ _2096_ _2110_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_119_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3648_ _1244_ _1245_ _1246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_20_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6436_ _0309_ clknet_leaf_98_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[3\]\[22\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_136_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6367_ _0240_ clknet_leaf_21_wb_clk_i soc.rom_encoder_0.input_buffer\[1\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3579_ _1163_ _1165_ _1177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_115_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5318_ soc.ram_encoder_0.data_out\[4\] _2551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_103_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6298_ _0173_ clknet_leaf_97_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[4\]\[27\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5249_ soc.ram_encoder_0.input_bits_left\[4\] _2497_ _2500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_102_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_2_wb_clk_i clknet_4_0_0_wb_clk_i clknet_leaf_2_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_72_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_141_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_117_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4620_ _2064_ _0151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_30_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_72_wb_clk_i clknet_4_15_0_wb_clk_i clknet_leaf_72_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_4551_ soc.spi_video_ram_1.fifo_in_data\[2\] soc.spi_video_ram_1.write_fifo.fifo_mem\[7\]\[2\]
+ _2023_ _2028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_144_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3502_ _1088_ _1089_ _1085_ _1102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4482_ soc.video_generator_1.v_count\[1\] _1980_ _1986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_144_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3433_ _0972_ _1029_ _1032_ _1037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_6221_ _0096_ clknet_leaf_140_wb_clk_i soc.video_generator_1.v_count\[5\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_143_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6152_ _0032_ clknet_leaf_61_wb_clk_i soc.ram_encoder_0.output_buffer\[13\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3364_ _0884_ _0970_ _0971_ _0879_ soc.cpu.PC.in\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5103_ soc.rom_encoder_0.initializing_step\[4\] soc.rom_encoder_0.initializing_step\[1\]
+ _1438_ _2384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_44_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3295_ _0849_ _0905_ _0906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_6083_ _3036_ _0643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5034_ net60 _2330_ _2346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_57_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5936_ soc.spi_video_ram_1.write_fifo.fifo_mem\[0\]\[4\] soc.spi_video_ram_1.fifo_in_data\[4\]
+ _2953_ _2958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5867_ _2915_ _0548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5798_ soc.cpu.PC.in\[6\] _2847_ _2861_ _2868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4818_ _2196_ _0218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_135_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4749_ soc.rom_encoder_0.request_data_out\[4\] _1481_ _2146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_123_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6419_ _0292_ clknet_leaf_129_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[3\]\[5\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xoutput58 net58 io_out[10] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput47 net47 io_oeb[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_89_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput69 net69 io_out[21] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_103_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3080_ soc.spi_video_ram_1.write_fifo.write_pointer\[2\] _0700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_94_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_36_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3982_ soc.ram_encoder_0.output_buffer\[9\] _1520_ _1530_ soc.ram_encoder_0.request_data_out\[5\]
+ _1546_ _1547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_6770_ _0612_ clknet_leaf_74_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[1\]\[12\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_51_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_0 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_94_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_62_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5721_ _2814_ _0503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5652_ soc.rom_loader.wait_fall_clk soc.rom_loader.rom_request _0175_ _2776_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_30_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5583_ soc.spi_video_ram_1.fifo_in_address\[7\] soc.spi_video_ram_1.write_fifo.fifo_mem\[5\]\[23\]
+ _2719_ _2732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_30_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4603_ _2054_ _0144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4534_ soc.spi_video_ram_1.fifo_in_data\[12\] _2007_ _2017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_117_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_144_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4465_ soc.spi_video_ram_1.state_counter\[7\] _1971_ _1974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3416_ _1018_ _1019_ _1020_ _1021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_6204_ _0007_ clknet_leaf_141_wb_clk_i soc.spi_video_ram_1.current_state\[4\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_4396_ _1609_ _1917_ _1918_ _1919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_112_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3347_ _0954_ _0955_ _0956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6135_ _0015_ clknet_leaf_2_wb_clk_i soc.video_generator_1.h_count\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_86_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6066_ _3027_ _0635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_58_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5017_ soc.ram_encoder_0.initializing_step\[4\] soc.ram_encoder_0.initializing_step\[3\]
+ _2331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3278_ net38 _0890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_27_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1806 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1839 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1817 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1828 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5919_ net16 _2947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_22_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_108_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_60_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_33_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4250_ soc.spi_video_ram_1.write_fifo.fifo_mem\[1\]\[8\] _1781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_141_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4181_ _1717_ _1718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3201_ _0758_ _0810_ _0815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_3132_ _0740_ _0743_ _0744_ _0746_ _0747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_95_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3063_ _0682_ _0683_ _0684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_36_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6822_ _0664_ clknet_leaf_54_wb_clk_i soc.ram_encoder_0.data_out\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_90_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3965_ soc.ram_encoder_0.request_address\[8\] _1513_ _1534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_6753_ _0595_ clknet_leaf_107_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[0\]\[24\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_32_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6684_ _0526_ net85 soc.cpu.PC.REG.data\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5704_ _2805_ _0495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3896_ _1132_ _1470_ _1472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5635_ soc.rom_loader.current_address\[9\] _2763_ _2765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_5566_ _1889_ _2707_ _2723_ _0439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5497_ _1488_ _2595_ _2678_ soc.ram_encoder_0.initializing_step\[2\] _0675_ _2679_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_4517_ _0009_ _0942_ _2008_ _0104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_137_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4448_ _1961_ _1962_ _0081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_144_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_120_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_59_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4379_ _1761_ _1902_ _1903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6118_ _0958_ _2897_ _3052_ _2551_ _0662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_100_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_86_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6049_ _3017_ _0628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_39_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_2_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_139_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_129_wb_clk_i clknet_4_3_0_wb_clk_i clknet_leaf_129_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_135_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_72_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_14_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3750_ _1345_ _1346_ _1218_ _1347_ _1138_ _1348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_3681_ _1272_ _1279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_127_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5420_ _2604_ _2620_ _2621_ _2622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_9_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5351_ _2572_ _2538_ _2573_ _0374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_57_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5282_ _2522_ _2504_ _2523_ _0355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_114_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4302_ _1702_ _1826_ _1829_ _1830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_114_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4233_ _0729_ _1765_ _1578_ _1692_ _1766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_68_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4164_ _1579_ _1702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_83_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4095_ _1645_ _1646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3115_ _0729_ _0732_ _0733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_70_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6805_ _0647_ clknet_leaf_82_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[2\]\[18\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_12_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4997_ _2316_ soc.rom_encoder_0.request_address\[9\] _2271_ _2317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_23_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6736_ _0578_ clknet_leaf_120_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[0\]\[7\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3948_ soc.ram_encoder_0.request_address\[4\] _1514_ _1520_ soc.ram_encoder_0.output_buffer\[1\]
+ _1521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_104_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_3879_ _1461_ _1268_ _1281_ _0014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_6667_ _0509_ clknet_leaf_118_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[6\]\[19\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5618_ _2746_ _2752_ _2753_ _0460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_6598_ net36 clknet_leaf_143_wb_clk_i soc.rom_encoder_0.data_out\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_117_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5549_ _2714_ _0431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_133_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_87_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_74_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2101 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2134 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2123 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2112 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2156 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2167 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2145 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2178 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_6_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_97_wb_clk_i clknet_4_11_0_wb_clk_i clknet_leaf_97_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_93_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_26_wb_clk_i clknet_4_5_0_wb_clk_i clknet_leaf_26_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_77_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4920_ soc.rom_encoder_0.input_buffer\[7\] _2241_ _2250_ _2267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_52_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4851_ soc.spi_video_ram_1.write_fifo.write_pointer\[2\] _0738_ _2216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_3802_ _1383_ _1390_ _1391_ _1392_ _1393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_4782_ soc.rom_encoder_0.output_buffer\[15\] _1417_ _1442_ soc.rom_encoder_0.request_data_out\[11\]
+ _2172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6521_ _0394_ clknet_leaf_57_wb_clk_i soc.ram_data_out\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3733_ soc.video_generator_1.v_count\[3\] _1129_ _1331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6452_ _0325_ clknet_leaf_51_wb_clk_i soc.cpu.ALU.ny vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3664_ soc.video_generator_1.h_count\[1\] soc.video_generator_1.h_count\[2\] _1215_
+ _1262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_5403_ net1 _2488_ _2608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6383_ _0256_ clknet_leaf_32_wb_clk_i soc.rom_encoder_0.request_data_out\[4\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3595_ _1133_ _1192_ _1193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_115_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5334_ soc.ram_encoder_0.request_data_out\[9\] _2545_ _2562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_142_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5265_ soc.ram_encoder_0.input_buffer\[3\] _2512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_87_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_134_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5196_ _2458_ _2269_ _1403_ _2459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4216_ _1594_ _1748_ _1749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_56_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4147_ _1611_ _1686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_84_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4078_ soc.spi_video_ram_1.output_buffer\[2\] _1612_ _1633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_71_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6719_ _0561_ clknet_leaf_8_wb_clk_i soc.hack_wait_clocks\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_7_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_59_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_144_wb_clk_i clknet_4_0_0_wb_clk_i clknet_leaf_144_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_42_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xcaravel_hack_soc_160 la_data_out[32] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xcaravel_hack_soc_171 la_data_out[43] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xcaravel_hack_soc_182 la_data_out[54] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_3380_ _0875_ _0986_ _0987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xcaravel_hack_soc_193 wbs_dat_o[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_69_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5050_ _2354_ _0292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4001_ _1562_ _0035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_111_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_1_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_81_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5952_ _2966_ _0582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4903_ _2254_ _2242_ _2255_ _0244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_18_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5883_ _2923_ _0556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4834_ _2204_ _0226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4765_ _1437_ _1482_ soc.rom_encoder_0.output_buffer\[12\] _2158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_14_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6504_ _0377_ clknet_leaf_65_wb_clk_i soc.ram_encoder_0.request_address\[1\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3716_ _1272_ _1313_ _1263_ _1314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4696_ _2108_ _2109_ _0182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6435_ _0308_ clknet_leaf_92_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[3\]\[21\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3647_ _1171_ _1180_ _1183_ _1245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_6366_ _0239_ clknet_leaf_21_wb_clk_i soc.rom_encoder_0.input_buffer\[0\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3578_ _1154_ _1172_ _1166_ _1175_ _1176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_143_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5317_ _2549_ _2542_ _2550_ _0363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_102_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6297_ _0172_ clknet_leaf_101_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[4\]\[26\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_130_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5248_ _2497_ _2498_ _2499_ _0345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_57_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5179_ _2436_ _2445_ _0330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_60_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_43_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_4_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_16_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_30_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_129_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4550_ _1708_ _2025_ _2027_ _0118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_7_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_143_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3501_ _1094_ _1087_ _1100_ _1101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_4481_ _1980_ _1984_ _1985_ _0091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_143_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_116_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3432_ _1026_ _1027_ _1034_ _1036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_6220_ _0095_ clknet_leaf_142_wb_clk_i soc.video_generator_1.v_count\[4\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_125_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_41_wb_clk_i clknet_4_7_0_wb_clk_i clknet_leaf_41_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_6151_ _0031_ clknet_leaf_62_wb_clk_i soc.ram_encoder_0.output_buffer\[12\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3363_ _0846_ soc.cpu.AReg.data\[5\] _0971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_83_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5102_ soc.rom_encoder_0.initializing_step\[2\] _2383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3294_ _0904_ soc.cpu.ALU.x\[2\] _0905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_44_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6082_ soc.spi_video_ram_1.write_fifo.fifo_mem\[2\]\[14\] soc.spi_video_ram_1.fifo_in_data\[14\]
+ _3031_ _3036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5033_ soc.ram_encoder_0.output_buffer\[18\] _1555_ _1529_ soc.ram_encoder_0.request_data_out\[14\]
+ _1559_ _2345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_66_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5935_ _2957_ _0574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5866_ soc.ram_encoder_0.address\[11\] soc.cpu.AReg.data\[11\] _2902_ _2915_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_22_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4817_ soc.spi_video_ram_1.fifo_in_address\[3\] soc.cpu.AReg.data\[3\] _2018_ _2196_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_21_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5797_ soc.cpu.PC.REG.data\[6\] _2866_ _2867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_22_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4748_ _2122_ _2144_ _2145_ _0199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_119_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4679_ soc.spi_video_ram_1.state_sram_clk_counter\[1\] _2095_ _2098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_116_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6418_ _0291_ clknet_leaf_9_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[3\]\[4\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_122_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput48 net48 io_oeb[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput59 net59 io_out[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_88_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6349_ _0223_ clknet_leaf_76_wb_clk_i soc.spi_video_ram_1.fifo_in_address\[8\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_131_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_103_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3981_ soc.ram_encoder_0.request_address\[12\] _1513_ _1546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_62_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_1 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_16_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5720_ soc.spi_video_ram_1.write_fifo.fifo_mem\[6\]\[13\] soc.spi_video_ram_1.fifo_in_data\[13\]
+ _2810_ _2814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_31_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5651_ net45 _2775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_50_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5582_ _2731_ _0447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4602_ soc.spi_video_ram_1.fifo_in_address\[11\] soc.spi_video_ram_1.write_fifo.fifo_mem\[7\]\[27\]
+ _2037_ _2054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_144_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4533_ _2003_ _1069_ _2016_ _0112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_144_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4464_ soc.spi_video_ram_1.state_counter\[7\] _1971_ _1973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_6203_ _0006_ clknet_leaf_135_wb_clk_i soc.spi_video_ram_1.current_state\[3\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_3415_ _1016_ _1020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4395_ _1144_ _1695_ _1918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_98_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3346_ _0947_ _0951_ _0955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6134_ _0014_ clknet_4_0_0_wb_clk_i soc.video_generator_1.h_count\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_113_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_100_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6065_ soc.spi_video_ram_1.write_fifo.fifo_mem\[2\]\[6\] soc.spi_video_ram_1.fifo_in_data\[6\]
+ _3020_ _3027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5016_ _1492_ _1508_ _2330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_3277_ _0887_ _0888_ _0889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_85_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1807 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1818 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1829 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5918_ _2945_ _2943_ _2946_ _0568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_107_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5849_ _0908_ _2903_ _2906_ _0539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_10_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4180_ soc.spi_video_ram_1.write_fifo.fifo_mem\[4\]\[2\] soc.spi_video_ram_1.write_fifo.fifo_mem\[5\]\[2\]
+ soc.spi_video_ram_1.write_fifo.fifo_mem\[6\]\[2\] soc.spi_video_ram_1.write_fifo.fifo_mem\[7\]\[2\]
+ _1593_ _1587_ _1717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_3200_ soc.spi_video_ram_1.output_buffer\[14\] soc.spi_video_ram_1.output_buffer\[15\]
+ _0783_ _0814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3131_ net87 soc.hack_clk_strobe soc.cpu.AReg.data\[14\] _0745_ _0746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_79_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_67_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3062_ soc.spi_video_ram_1.state_sram_clk_counter\[3\] soc.spi_video_ram_1.state_sram_clk_counter\[2\]
+ _0683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_82_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6821_ _0663_ clknet_leaf_54_wb_clk_i soc.ram_encoder_0.data_out\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_63_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3964_ _1510_ _1532_ _1533_ _0027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_51_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6752_ _0594_ clknet_leaf_103_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[0\]\[23\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6683_ _0525_ net84 soc.cpu.PC.REG.data\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5703_ soc.spi_video_ram_1.write_fifo.fifo_mem\[6\]\[5\] soc.spi_video_ram_1.fifo_in_data\[5\]
+ _2799_ _2805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3895_ _1132_ _1470_ _1471_ _0020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5634_ soc.rom_loader.current_address\[9\] _2763_ _2764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_31_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5565_ soc.spi_video_ram_1.fifo_in_data\[14\] _2708_ _2723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5496_ soc.ram_encoder_0.initializing_step\[1\] soc.ram_encoder_0.initializing_step\[0\]
+ _2597_ _2678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_105_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4516_ soc.spi_video_ram_1.fifo_in_data\[3\] _2007_ _2008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4447_ soc.spi_video_ram_1.state_counter\[1\] soc.spi_video_ram_1.state_counter\[0\]
+ _1962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_113_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6117_ _0942_ _2897_ _3052_ _2549_ _0661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_98_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4378_ _1901_ _1902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3329_ _0925_ _0935_ _0939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_74_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6048_ soc.spi_video_ram_1.fifo_in_address\[12\] soc.spi_video_ram_1.write_fifo.fifo_mem\[1\]\[28\]
+ _2985_ _3017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_2316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_4_8_0_wb_clk_i clknet_0_wb_clk_i clknet_4_8_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_42_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_40_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_32_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3680_ _1217_ _1218_ _1278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_40_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5350_ soc.ram_encoder_0.request_data_out\[14\] _2566_ _2573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5281_ soc.ram_encoder_0.input_buffer\[4\] _2503_ _2508_ _2523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4301_ _1761_ _1828_ _1829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_5_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4232_ _1693_ _1694_ _1765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4163_ soc.spi_video_ram_1.write_fifo.fifo_mem\[2\]\[1\] soc.spi_video_ram_1.write_fifo.fifo_mem\[3\]\[1\]
+ _1600_ _1701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_67_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4094_ _0674_ _1427_ _1424_ _1645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_3114_ soc.spi_video_ram_1.state_sram_clk_counter\[6\] _0715_ _0717_ _0731_ _0732_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__or4_1
XFILLER_110_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_51_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4996_ soc.cpu.PC.REG.data\[9\] soc.rom_loader.current_address\[9\] _2292_ _2316_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6804_ _0646_ clknet_leaf_84_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[2\]\[17\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_24_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3947_ _1519_ _1520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_6735_ _0577_ clknet_leaf_124_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[0\]\[6\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_17_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6666_ _0508_ clknet_leaf_84_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[6\]\[18\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_31_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3878_ _0689_ _1461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_5617_ soc.rom_loader.current_address\[3\] _2751_ _2753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_6597_ net35 clknet_leaf_94_wb_clk_i soc.rom_encoder_0.data_out\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5548_ soc.spi_video_ram_1.fifo_in_data\[6\] soc.spi_video_ram_1.write_fifo.fifo_mem\[5\]\[6\]
+ _2705_ _2714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_132_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_117_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5479_ _1955_ _2542_ _2666_ _0409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_101_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2135 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2124 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2113 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2102 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2157 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2168 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2146 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_15_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2179 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_66_wb_clk_i clknet_4_13_0_wb_clk_i clknet_leaf_66_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_80_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_61_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4850_ _0694_ _2213_ _2215_ _0231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3801_ _0761_ _0766_ _1383_ _1392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_1990 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6520_ _0393_ clknet_leaf_47_wb_clk_i soc.ram_data_out\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4781_ _1671_ _2170_ _2171_ _0206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_20_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3732_ _1190_ _1131_ _1327_ _1329_ _1330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_6451_ _0324_ clknet_leaf_51_wb_clk_i soc.cpu.ALU.f vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_9_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3663_ _1260_ _1261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_5402_ soc.ram_encoder_0.request_data_out\[0\] _2606_ _2607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6382_ _0255_ clknet_leaf_11_wb_clk_i soc.rom_encoder_0.request_data_out\[3\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_114_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5333_ soc.ram_encoder_0.data_out\[9\] _2561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_86_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3594_ _1189_ _1191_ _1192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_88_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5264_ _2510_ _2504_ _2511_ _0349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5195_ _1407_ _2224_ _2458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4215_ soc.spi_video_ram_1.write_fifo.fifo_mem\[3\]\[6\] _1748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_68_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4146_ soc.spi_video_ram_1.output_buffer\[23\] _1685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_29_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4077_ _1581_ _1624_ _1631_ _1609_ _1632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_43_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4979_ soc.cpu.PC.REG.data\[4\] soc.rom_loader.current_address\[4\] _2292_ _2304_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_133_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6718_ _0560_ clknet_leaf_50_wb_clk_i soc.rom_encoder_0.write_enable vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_109_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6649_ _0491_ clknet_leaf_125_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[6\]\[1\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_125_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_129_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_109_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xcaravel_hack_soc_150 la_data_out[21] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xclkbuf_leaf_113_wb_clk_i clknet_4_8_0_wb_clk_i clknet_leaf_113_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
Xcaravel_hack_soc_183 la_data_out[55] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xcaravel_hack_soc_161 la_data_out[33] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xcaravel_hack_soc_172 la_data_out[44] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_112_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xcaravel_hack_soc_194 wbs_dat_o[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_85_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4000_ _1561_ soc.ram_encoder_0.output_buffer\[16\] _1509_ _1562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_111_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_38_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_19_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5951_ soc.spi_video_ram_1.write_fifo.fifo_mem\[0\]\[11\] soc.spi_video_ram_1.fifo_in_data\[11\]
+ _2964_ _2966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_52_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4902_ soc.rom_encoder_0.input_buffer\[1\] _2243_ _2250_ _2255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_33_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5882_ soc.boot_loading_offset\[1\] _2921_ _2922_ _2923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4833_ soc.spi_video_ram_1.fifo_in_address\[11\] soc.cpu.AReg.data\[11\] _0748_ _2204_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_21_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4764_ _2122_ _2156_ _2157_ _0203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_119_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6503_ _0376_ clknet_leaf_64_wb_clk_i soc.ram_encoder_0.request_address\[0\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3715_ _1261_ _1312_ _1239_ _1313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_101_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4695_ soc.spi_video_ram_1.state_sram_clk_counter\[6\] _2106_ _2096_ _2109_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6434_ _0307_ clknet_leaf_118_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[3\]\[20\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3646_ _1242_ _1243_ _1244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_115_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6365_ _0238_ clknet_leaf_3_wb_clk_i soc.rom_encoder_0.input_bits_left\[4\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3577_ _1173_ _1156_ _1171_ _1174_ _1175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XFILLER_142_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5316_ soc.ram_encoder_0.request_data_out\[3\] _2545_ _2550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_88_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6296_ _0171_ clknet_leaf_105_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[4\]\[25\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5247_ soc.ram_encoder_0.input_bits_left\[3\] _2495_ _2499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_103_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5178_ soc.cpu.instruction\[13\] _2393_ _2444_ _2445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_69_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4129_ _1674_ _0050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_72_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_24_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3500_ _1096_ _1099_ _1100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4480_ soc.video_generator_1.v_count\[0\] _1458_ _1985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_144_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3431_ _1026_ _1027_ _1034_ _1035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_124_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6150_ _0030_ clknet_leaf_61_wb_clk_i soc.ram_encoder_0.output_buffer\[11\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_98_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3362_ _0922_ _0960_ _0969_ _0970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XTAP_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5101_ _2380_ _2381_ _1438_ _2382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_32_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3293_ _0850_ _0904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_6081_ _3035_ _0642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xclkbuf_4_10_0_wb_clk_i clknet_0_wb_clk_i clknet_4_10_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XTAP_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5032_ _2330_ _2343_ _2344_ _0676_ _0284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
Xclkbuf_leaf_81_wb_clk_i clknet_4_14_0_wb_clk_i clknet_leaf_81_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_57_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_10_wb_clk_i clknet_4_1_0_wb_clk_i clknet_leaf_10_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_81_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5934_ soc.spi_video_ram_1.write_fifo.fifo_mem\[0\]\[3\] soc.spi_video_ram_1.fifo_in_data\[3\]
+ _2953_ _2957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5865_ _2914_ _0547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4816_ _2195_ _0217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_21_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5796_ soc.cpu.PC.REG.data\[5\] _2863_ _2866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_22_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4747_ soc.rom_encoder_0.output_buffer\[11\] _2138_ _2145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4678_ _2095_ _2097_ _0176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3629_ _1198_ _1226_ _1227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6417_ _0290_ clknet_leaf_9_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[3\]\[3\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6348_ _0222_ clknet_4_15_0_wb_clk_i soc.spi_video_ram_1.fifo_in_address\[7\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
Xoutput49 net49 io_oeb[13] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_103_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6279_ _0154_ clknet_leaf_121_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[4\]\[8\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_102_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_40_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_126_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3980_ _1510_ _1544_ _1545_ _0031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_50_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5650_ _2746_ _2774_ _0471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4601_ _2053_ _0143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_129_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5581_ soc.spi_video_ram_1.fifo_in_address\[6\] soc.spi_video_ram_1.write_fifo.fifo_mem\[5\]\[22\]
+ _2719_ _2731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4532_ soc.spi_video_ram_1.fifo_in_data\[11\] _2007_ _2016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_11_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_7_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4463_ _1961_ _1971_ _1972_ _0086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_3414_ _1000_ _1006_ _1007_ _1019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_6202_ _0005_ clknet_leaf_137_wb_clk_i soc.spi_video_ram_1.current_state\[2\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_125_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4394_ _1913_ _1914_ _1915_ _1916_ _1591_ _1761_ _1917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_112_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3345_ soc.cpu.ALU.f _0954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6133_ _0013_ clknet_leaf_2_wb_clk_i soc.display_clks_before_active\[0\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_112_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3276_ soc.ram_data_out\[1\] _0869_ _0888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_86_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6064_ _3026_ _0634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5015_ _2329_ _0282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1819 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1808 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5917_ soc.gpio_i_stored\[1\] _2943_ _2531_ _2946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_41_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5848_ soc.ram_encoder_0.address\[2\] _2903_ _2906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_21_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5779_ soc.cpu.PC.REG.data\[0\] soc.cpu.PC.REG.data\[1\] _2853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_108_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_104_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_29_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3130_ soc.cpu.AReg.data\[13\] _0745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_68_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3061_ soc.spi_video_ram_1.state_sram_clk_counter\[7\] soc.spi_video_ram_1.state_sram_clk_counter\[6\]
+ soc.spi_video_ram_1.state_sram_clk_counter\[5\] soc.spi_video_ram_1.state_sram_clk_counter\[4\]
+ _0682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_48_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6820_ _0662_ clknet_leaf_54_wb_clk_i soc.ram_encoder_0.data_out\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_91_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3963_ soc.ram_encoder_0.output_buffer\[8\] _1527_ _1533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6751_ _0593_ clknet_leaf_97_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[0\]\[22\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6682_ _0524_ net84 soc.cpu.PC.REG.data\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5702_ _2804_ _0494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_32_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3894_ _1132_ _1470_ _1462_ _1471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5633_ _2746_ _2762_ _2763_ _0465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_5564_ _1866_ _2707_ _2722_ _0438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4515_ _0748_ _2007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_144_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5495_ _1516_ _2676_ _2677_ _2471_ _0414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_4446_ soc.spi_video_ram_1.state_counter\[0\] _1961_ _0080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_101_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4377_ soc.spi_video_ram_1.write_fifo.fifo_mem\[4\]\[15\] soc.spi_video_ram_1.write_fifo.fifo_mem\[5\]\[15\]
+ soc.spi_video_ram_1.write_fifo.fifo_mem\[6\]\[15\] soc.spi_video_ram_1.write_fifo.fifo_mem\[7\]\[15\]
+ _1583_ _1586_ _1901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_113_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6116_ _0920_ _2897_ _3052_ _2547_ _0660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_3328_ _0925_ _0935_ _0937_ _0938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XTAP_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3259_ soc.gpio_i_stored\[0\] _0867_ _0868_ net29 _0871_ _0872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_85_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_74_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_27_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6047_ _3016_ _0627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_138_wb_clk_i clknet_4_2_0_wb_clk_i clknet_leaf_138_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_58_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_18_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5280_ soc.ram_encoder_0.input_buffer\[8\] _2522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4300_ _1827_ _1828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4231_ _1753_ _1763_ _0703_ _1608_ _1764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_142_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4162_ _1595_ soc.spi_video_ram_1.write_fifo.fifo_mem\[0\]\[1\] _1699_ _1700_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4093_ _1643_ _1644_ _0044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_68_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_56_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3113_ soc.spi_video_ram_1.state_sram_clk_counter\[7\] _0730_ _0731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_55_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_64_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4995_ _2315_ _0276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6803_ _0645_ clknet_leaf_80_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[2\]\[16\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_23_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3946_ _1515_ _1516_ _1518_ _1519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_51_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6734_ _0576_ clknet_leaf_128_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[0\]\[5\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_136_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6665_ _0507_ clknet_leaf_86_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[6\]\[17\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_20_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3877_ _1216_ _1460_ _0013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6596_ net34 clknet_leaf_41_wb_clk_i soc.rom_encoder_0.data_out\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5616_ soc.rom_loader.current_address\[3\] _2751_ _2752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_118_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5547_ _1740_ _2707_ _2713_ _0430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_3_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5478_ _2492_ _2535_ soc.ram_encoder_0.sram_sio_oe _2666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_144_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4429_ _1578_ _1947_ _1948_ _0076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_87_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2125 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2114 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2103 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2158 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2147 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2136 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2169 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_14_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout84 net86 net84 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_7_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_108_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_124_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_96_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4780_ soc.rom_encoder_0.output_buffer\[18\] _2138_ _2171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3800_ _0758_ soc.spi_video_ram_1.output_buffer\[1\] _0775_ _1391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_33_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1991 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1980 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3731_ soc.video_generator_1.h_count\[4\] _1328_ _1329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_118_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_35_wb_clk_i clknet_4_7_0_wb_clk_i clknet_leaf_35_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_6450_ _0323_ clknet_leaf_51_wb_clk_i soc.cpu.ALU.no vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3662_ _1247_ _1256_ _1259_ _1260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_5401_ _2605_ _2606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_62_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6381_ _0254_ clknet_leaf_11_wb_clk_i soc.rom_encoder_0.request_data_out\[2\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3593_ _1190_ _1132_ _1131_ _1191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_5332_ _2559_ _2542_ _2560_ _0368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_141_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5263_ net3 _2505_ _2508_ _2511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_102_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5194_ _2457_ _0333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4214_ _0801_ _1686_ _1697_ _1747_ _0062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4145_ _1522_ _1683_ _1684_ _0056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_69_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_29_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4076_ _1592_ _1627_ _1630_ _1605_ _1631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_37_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_51_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4978_ _2272_ _2302_ _2303_ _0271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_52_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3929_ soc.ram_encoder_0.current_state\[0\] _1502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_20_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6717_ _0559_ clknet_leaf_8_wb_clk_i soc.boot_loading_offset\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_137_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6648_ _0490_ clknet_leaf_12_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[6\]\[0\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_50_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_30_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6579_ _0452_ clknet_4_10_0_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[5\]\[27\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_121_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_10_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xcaravel_hack_soc_140 la_data_out[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xcaravel_hack_soc_184 la_data_out[56] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xcaravel_hack_soc_173 la_data_out[45] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xcaravel_hack_soc_162 la_data_out[34] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xcaravel_hack_soc_151 la_data_out[22] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_123_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xcaravel_hack_soc_195 wbs_dat_o[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_112_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5950_ _2965_ _0581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_53_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4901_ soc.rom_encoder_0.input_buffer\[5\] _2254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5881_ soc.boot_loading_offset\[1\] _2921_ _0689_ _2922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4832_ _2203_ _0225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_60_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4763_ soc.rom_encoder_0.output_buffer\[15\] _2138_ _2157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_53_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6502_ _0375_ clknet_leaf_46_wb_clk_i soc.ram_encoder_0.request_data_out\[15\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4694_ soc.spi_video_ram_1.state_sram_clk_counter\[6\] _2106_ _2108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_3714_ _1286_ _1269_ _1301_ _1312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_135_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6433_ _0306_ clknet_leaf_89_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[3\]\[19\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_106_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3645_ _1167_ _1163_ _1243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_115_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6364_ _0237_ clknet_leaf_3_wb_clk_i soc.rom_encoder_0.input_bits_left\[3\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3576_ soc.boot_loading_offset\[2\] _1156_ _1147_ _1174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_143_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5315_ soc.ram_encoder_0.data_out\[3\] _2549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_88_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6295_ _0170_ clknet_leaf_106_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[4\]\[24\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5246_ _2488_ _2494_ _2498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_69_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5177_ _2262_ _2413_ _2414_ _2443_ _2444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_68_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4128_ soc.rom_encoder_0.output_buffer\[3\] _1671_ _1672_ soc.rom_encoder_0.request_address\[2\]
+ _1674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_72_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4059_ soc.spi_video_ram_1.write_fifo.fifo_mem\[5\]\[18\] _1615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_83_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_16_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_35_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3430_ _1033_ _1034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3361_ _0954_ _0967_ _0968_ _0969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_124_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5100_ _2221_ _1425_ _2381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_3_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6080_ soc.spi_video_ram_1.write_fifo.fifo_mem\[2\]\[13\] soc.spi_video_ram_1.fifo_in_data\[13\]
+ _3031_ _3035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5031_ net59 _2330_ _2344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_111_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_98_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3292_ _0884_ _0902_ _0903_ soc.cpu.PC.in\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_38_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_50_wb_clk_i clknet_4_6_0_wb_clk_i clknet_leaf_50_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_81_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_34_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5933_ _2956_ _0573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5864_ soc.ram_encoder_0.address\[10\] soc.cpu.AReg.data\[10\] _2902_ _2914_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_90_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4815_ soc.spi_video_ram_1.fifo_in_address\[2\] soc.cpu.AReg.data\[2\] _2018_ _2195_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_21_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5795_ _2846_ _2864_ _2865_ _0525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_21_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4746_ soc.rom_encoder_0.request_address\[10\] _1650_ _2125_ soc.rom_encoder_0.output_buffer\[7\]
+ _2143_ _2144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_107_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4677_ soc.spi_video_ram_1.state_sram_clk_counter\[0\] _2094_ _2096_ _2097_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_134_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6416_ _0289_ clknet_leaf_10_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[3\]\[2\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3628_ _1190_ _1135_ _1197_ _1226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6347_ _0221_ clknet_leaf_75_wb_clk_i soc.spi_video_ram_1.fifo_in_address\[6\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3559_ soc.boot_loading_offset\[2\] _1156_ _1157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_103_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6278_ _0153_ clknet_leaf_125_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[4\]\[7\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_76_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5229_ _2476_ _2482_ _2484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_57_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_53_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_80_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_3 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_16_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4600_ soc.spi_video_ram_1.fifo_in_address\[10\] soc.spi_video_ram_1.write_fifo.fifo_mem\[7\]\[26\]
+ _2037_ _2053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5580_ _2730_ _0446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_117_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4531_ _2003_ _1058_ _2015_ _0111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4462_ soc.spi_video_ram_1.state_counter\[6\] _1969_ _1972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_144_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3413_ _0945_ _0981_ _1004_ _1018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_6201_ _0004_ clknet_leaf_133_wb_clk_i soc.spi_video_ram_1.current_state\[1\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_113_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4393_ soc.spi_video_ram_1.write_fifo.fifo_mem\[6\]\[22\] soc.spi_video_ram_1.write_fifo.fifo_mem\[7\]\[22\]
+ _1584_ _1916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_140_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3344_ _0945_ _0952_ _0953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6132_ _0012_ clknet_leaf_1_wb_clk_i net67 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3275_ soc.cpu.instruction\[12\] _0887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XTAP_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6063_ soc.spi_video_ram_1.write_fifo.fifo_mem\[2\]\[5\] soc.spi_video_ram_1.fifo_in_data\[5\]
+ _3020_ _3026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_85_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5014_ _2328_ soc.rom_encoder_0.request_address\[14\] _2271_ _2329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5916_ net15 _2945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_81_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5847_ _2905_ _0538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_22_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5778_ _2846_ _2850_ _2852_ _2849_ _0521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_4729_ soc.rom_encoder_0.output_buffer\[7\] _1670_ _2131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_135_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_8_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3060_ soc.spi_video_ram_1.state_sram_clk_counter\[1\] _0681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_82_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_17_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6750_ _0592_ clknet_leaf_97_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[0\]\[21\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3962_ soc.ram_encoder_0.output_buffer\[4\] _1520_ _1530_ soc.ram_encoder_0.request_data_out\[0\]
+ _1531_ _1532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_92_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5701_ soc.spi_video_ram_1.write_fifo.fifo_mem\[6\]\[4\] soc.spi_video_ram_1.fifo_in_data\[4\]
+ _2799_ _2804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_32_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6681_ _0523_ net84 soc.cpu.PC.REG.data\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_50_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3893_ _1460_ _1469_ _1470_ _0019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_5632_ soc.rom_loader.current_address\[8\] soc.rom_loader.current_address\[7\] _2759_
+ _2763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_129_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5563_ soc.spi_video_ram_1.fifo_in_data\[13\] _2708_ _2722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_117_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4514_ _0009_ _0920_ _2006_ _0103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_8_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5494_ soc.ram_encoder_0.initializing_step\[1\] _2598_ _2677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_137_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4445_ _1960_ _1961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_144_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4376_ soc.spi_video_ram_1.write_fifo.fifo_mem\[0\]\[15\] soc.spi_video_ram_1.write_fifo.fifo_mem\[1\]\[15\]
+ soc.spi_video_ram_1.write_fifo.fifo_mem\[2\]\[15\] soc.spi_video_ram_1.write_fifo.fifo_mem\[3\]\[15\]
+ _1724_ _1587_ _1900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_112_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6115_ _0902_ _2897_ _3052_ _2544_ _0659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_99_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_86_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3327_ _0917_ _0936_ _0916_ _0937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XTAP_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3258_ soc.cpu.instruction\[12\] _0870_ _0871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6046_ soc.spi_video_ram_1.fifo_in_address\[11\] soc.spi_video_ram_1.write_fifo.fifo_mem\[1\]\[27\]
+ _2985_ _3016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_2307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3189_ _0799_ _0800_ _0801_ _0802_ _0758_ _0776_ _0803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_2329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_14_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_120_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_131_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_2_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_107_wb_clk_i clknet_4_10_0_wb_clk_i clknet_leaf_107_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_32_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4230_ _0685_ _1762_ _1763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4161_ _1601_ _1698_ _1591_ _1699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_110_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4092_ soc.ram_encoder_0.output_bits_left\[2\] _1634_ _1644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3112_ soc.spi_video_ram_1.state_sram_clk_counter\[5\] soc.spi_video_ram_1.state_sram_clk_counter\[4\]
+ _0730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_83_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6802_ _0644_ clknet_leaf_73_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[2\]\[15\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4994_ _2314_ soc.rom_encoder_0.request_address\[8\] _2271_ _2315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_23_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3945_ _1504_ _1517_ _1518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_6733_ _0575_ clknet_leaf_130_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[0\]\[4\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6664_ _0506_ clknet_leaf_86_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[6\]\[16\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5615_ _2746_ _2750_ _2751_ _0459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_3876_ _1459_ _1460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6595_ net33 clknet_leaf_33_wb_clk_i soc.rom_encoder_0.data_out\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5546_ soc.spi_video_ram_1.fifo_in_data\[5\] _2708_ _2713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_144_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5477_ _2662_ _2664_ _2665_ _0408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_2_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4428_ soc.spi_video_ram_1.output_buffer\[4\] _1611_ _1948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_132_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4359_ _1593_ _1883_ _1590_ _1884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_74_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6029_ _3007_ _0618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xclkbuf_leaf_5_wb_clk_i clknet_4_1_0_wb_clk_i clknet_leaf_5_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_46_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2126 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2115 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2104 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2159 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2148 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2137 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout85 net86 net85 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_7_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_109_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_13_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_97_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1970 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1992 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1981 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3730_ _1132_ _1328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3661_ _1126_ _1257_ _1258_ _1259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5400_ _1493_ _1496_ _2605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
Xclkbuf_leaf_75_wb_clk_i clknet_4_15_0_wb_clk_i clknet_leaf_75_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_6380_ _0253_ clknet_leaf_25_wb_clk_i soc.rom_encoder_0.request_data_out\[1\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3592_ soc.video_generator_1.h_count\[5\] _1190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_5331_ soc.ram_encoder_0.request_data_out\[8\] _2545_ _2560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_86_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5262_ soc.ram_encoder_0.input_buffer\[2\] _2510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_114_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5193_ _1461_ _2456_ _2457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_4213_ _0685_ _1739_ _1746_ _1747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_4144_ soc.ram_encoder_0.output_buffer\[1\] _1509_ _1684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_56_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4075_ _1601_ soc.spi_video_ram_1.write_fifo.fifo_mem\[6\]\[17\] _1629_ _1591_ _1630_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_64_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4977_ soc.rom_encoder_0.request_address\[3\] _2272_ _2303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6716_ _0558_ clknet_leaf_9_wb_clk_i soc.boot_loading_offset\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_3928_ _1488_ _1500_ _1501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6647_ _0489_ net89 soc.cpu.ALU.x\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3859_ net65 _1432_ _1446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6578_ _0451_ clknet_leaf_103_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[5\]\[26\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_118_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5529_ soc.hack_clock_0.counter\[6\] _2701_ _2702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_106_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_42_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_7_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xcaravel_hack_soc_141 la_data_out[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xcaravel_hack_soc_130 la_data_out[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xcaravel_hack_soc_152 la_data_out[23] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xcaravel_hack_soc_174 la_data_out[46] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_108_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xcaravel_hack_soc_163 la_data_out[35] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xcaravel_hack_soc_185 la_data_out[57] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_124_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xcaravel_hack_soc_196 wbs_dat_o[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_2_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_122_wb_clk_i clknet_4_9_0_wb_clk_i clknet_leaf_122_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_19_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_37_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4900_ _2252_ _2242_ _2253_ _0243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_18_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5880_ _1461_ _2920_ _2921_ _0555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_4831_ soc.spi_video_ram_1.fifo_in_address\[10\] soc.cpu.AReg.data\[10\] _0748_ _2203_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_61_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4762_ soc.rom_encoder_0.request_address\[14\] _1650_ _2124_ soc.rom_encoder_0.output_buffer\[11\]
+ _2155_ _2156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_60_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6501_ _0374_ clknet_leaf_49_wb_clk_i soc.ram_encoder_0.request_data_out\[14\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4693_ _2106_ _2107_ _0181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_14_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3713_ _1276_ _1311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_128_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6432_ _0305_ clknet_leaf_82_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[3\]\[18\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3644_ _1127_ _1211_ _1242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_127_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6363_ _0236_ clknet_leaf_3_wb_clk_i soc.rom_encoder_0.input_bits_left\[2\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3575_ _1166_ _1169_ _1173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_143_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5314_ _2547_ _2542_ _2548_ _0362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6294_ _0169_ clknet_leaf_104_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[4\]\[23\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_143_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5245_ soc.ram_encoder_0.input_bits_left\[3\] _2495_ _2497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_88_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5176_ soc.rom_encoder_0.request_data_out\[13\] _2394_ _2443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_57_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4127_ _1673_ _0049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_84_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4058_ soc.spi_video_ram_1.write_fifo.fifo_mem\[0\]\[18\] soc.spi_video_ram_1.write_fifo.fifo_mem\[1\]\[18\]
+ soc.spi_video_ram_1.write_fifo.fifo_mem\[2\]\[18\] soc.spi_video_ram_1.write_fifo.fifo_mem\[3\]\[18\]
+ _1585_ _1588_ _1614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_24_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_143_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3360_ _0962_ _0966_ _0968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_125_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5030_ soc.ram_encoder_0.output_buffer\[17\] _1555_ _1529_ soc.ram_encoder_0.request_data_out\[13\]
+ _1559_ _2343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_97_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3291_ _0846_ soc.cpu.DMuxJMP.sel\[1\] soc.cpu.AReg.data\[1\] _0881_ _0903_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai22_1
XTAP_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5932_ soc.spi_video_ram_1.write_fifo.fifo_mem\[0\]\[2\] soc.spi_video_ram_1.fifo_in_data\[2\]
+ _2953_ _2956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_80_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5863_ _2913_ _0546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_61_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5794_ soc.cpu.PC.in\[5\] _2847_ _2861_ _2865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4814_ _2194_ _0216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_21_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4745_ soc.rom_encoder_0.request_data_out\[3\] _1481_ _2143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
Xclkbuf_leaf_90_wb_clk_i clknet_4_11_0_wb_clk_i clknet_leaf_90_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_21_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4676_ soc.spi_video_ram_1.current_state\[2\] net68 _2096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_116_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3627_ _1144_ _1173_ _1171_ _1224_ _1225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6415_ _0288_ clknet_leaf_129_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[3\]\[1\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_143_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6346_ _0220_ clknet_leaf_76_wb_clk_i soc.spi_video_ram_1.fifo_in_address\[5\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_3558_ _1149_ _1150_ _1156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_131_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3489_ _1088_ _1089_ _1085_ _0954_ _1090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_6277_ _0152_ clknet_leaf_123_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[4\]\[6\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5228_ _2480_ _2478_ _2481_ _2483_ _0690_ _0341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_5159_ soc.rom_encoder_0.request_data_out\[9\] _2394_ _2430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_71_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_122_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_138_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_21_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_4_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_31_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_43_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4530_ soc.spi_video_ram_1.fifo_in_data\[10\] _2007_ _2015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_7_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4461_ soc.spi_video_ram_1.state_counter\[6\] _1969_ _1971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_144_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3412_ _1005_ _1008_ _1016_ _1017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_6200_ _0003_ clknet_leaf_135_wb_clk_i soc.spi_video_ram_1.current_state\[0\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_98_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4392_ soc.spi_video_ram_1.write_fifo.fifo_mem\[4\]\[22\] soc.spi_video_ram_1.write_fifo.fifo_mem\[5\]\[22\]
+ _1584_ _1915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6131_ _0011_ clknet_leaf_8_wb_clk_i net66 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_98_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3343_ _0947_ _0951_ _0952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3274_ _0849_ _0885_ _0886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6062_ _3025_ _0633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5013_ soc.cpu.PC.REG.data\[14\] soc.rom_loader.current_address\[14\] _2292_ _2328_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_79_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5915_ _2941_ _2943_ _2944_ _0567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_53_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5846_ soc.ram_encoder_0.address\[1\] soc.cpu.AReg.data\[1\] _2903_ _2905_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_50_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_10_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5777_ soc.cpu.PC.in\[1\] _2851_ _2852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_22_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4728_ soc.rom_encoder_0.output_buffer\[3\] _2125_ _2130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_108_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4659_ _2084_ _0170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_89_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6329_ _0204_ clknet_leaf_4_wb_clk_i soc.rom_encoder_0.output_buffer\[16\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_103_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_91_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_29_wb_clk_i clknet_4_5_0_wb_clk_i clknet_leaf_29_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_63_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3961_ soc.ram_encoder_0.request_address\[7\] _1514_ _1531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_63_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5700_ _2803_ _0493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_50_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6680_ _0522_ net84 soc.cpu.PC.REG.data\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3892_ _1190_ _1131_ _1466_ _1470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_5631_ soc.rom_loader.current_address\[7\] _2759_ soc.rom_loader.current_address\[8\]
+ _2762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_85_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5562_ _2721_ _0437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4513_ soc.spi_video_ram_1.fifo_in_data\[2\] _2003_ _2006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5493_ _1488_ _2595_ _2676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_144_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_144_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4444_ _0709_ _1959_ _0674_ _1960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_98_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4375_ _1811_ _1898_ _1899_ _0071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6114_ _0878_ _2897_ _3052_ _2541_ _0658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_101_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3326_ _0906_ _0915_ _0936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6045_ _3015_ _0626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3257_ soc.ram_data_out\[0\] _0869_ _0870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3188_ soc.spi_video_ram_1.output_buffer\[16\] _0802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_2319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5829_ soc.cpu.PC.REG.data\[14\] _2890_ _2891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_22_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_17_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4160_ soc.spi_video_ram_1.write_fifo.fifo_mem\[1\]\[1\] _1698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_96_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3111_ soc.spi_video_ram_1.current_state\[4\] _0729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_4091_ soc.ram_encoder_0.output_bits_left\[2\] _1557_ _1634_ _1643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_110_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6801_ _0643_ clknet_leaf_99_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[2\]\[14\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4993_ soc.cpu.PC.REG.data\[8\] soc.rom_loader.current_address\[8\] _2292_ _2314_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_17_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3944_ _1500_ _1511_ _1517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6732_ _0574_ clknet_leaf_129_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[0\]\[3\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_143_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6663_ _0505_ clknet_leaf_93_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[6\]\[15\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_17_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3875_ net18 _1458_ _1459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_104_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5614_ soc.rom_loader.current_address\[2\] soc.rom_loader.current_address\[1\] _2744_
+ _2751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_6594_ net32 clknet_leaf_41_wb_clk_i soc.rom_encoder_0.data_out\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5545_ _2712_ _0429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_117_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5476_ net81 _2662_ _0690_ _2665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_133_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4427_ _1581_ _1939_ _1946_ _1609_ _1947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_63_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4358_ soc.spi_video_ram_1.write_fifo.fifo_mem\[1\]\[14\] _1883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_100_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3309_ soc.cpu.ALU.no _0919_ _0920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XTAP_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4289_ _1817_ _1818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_101_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6028_ soc.spi_video_ram_1.fifo_in_address\[2\] soc.spi_video_ram_1.write_fifo.fifo_mem\[1\]\[18\]
+ _2999_ _3007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_58_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2116 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2105 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2149 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2138 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2127 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout86 soc.cpu.AReg.clk net86 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyd_1
XFILLER_109_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_108_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_6_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_2_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1960 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1993 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1982 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1971 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3660_ _1127_ _1211_ _1243_ _1258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_127_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3591_ soc.video_generator_1.h_count\[8\] soc.video_generator_1.h_count\[9\] _1189_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_5330_ soc.ram_encoder_0.data_out\[8\] _2559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_6_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5261_ _2507_ _2504_ _2509_ _0348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xclkbuf_4_7_0_wb_clk_i clknet_0_wb_clk_i clknet_4_7_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_4212_ _1592_ _1742_ _1745_ _1605_ _1746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_48_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xclkbuf_leaf_44_wb_clk_i clknet_4_7_0_wb_clk_i clknet_leaf_44_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_96_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5192_ net62 _2453_ _2455_ _2456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4143_ soc.ram_encoder_0.request_address\[0\] _1514_ _1683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_95_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4074_ _1594_ _1628_ _1629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_28_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4976_ _2293_ soc.rom_loader.current_address\[3\] _2301_ _2302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_52_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6715_ _0557_ clknet_leaf_9_wb_clk_i soc.boot_loading_offset\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3927_ soc.ram_encoder_0.current_state\[2\] _1490_ _1500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6646_ _0488_ net90 soc.cpu.ALU.x\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3858_ soc.rom_encoder_0.output_buffer\[17\] _1436_ _1441_ _1444_ _1445_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_50_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6577_ _0450_ clknet_leaf_111_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[5\]\[25\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3789_ _0775_ _0790_ _1380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_30_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5528_ soc.hack_clock_0.counter\[5\] _2698_ _2701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5459_ soc.ram_data_out\[12\] _2604_ _2651_ _2652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_105_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xcaravel_hack_soc_120 io_out[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_136_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xcaravel_hack_soc_131 la_data_out[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xcaravel_hack_soc_142 la_data_out[13] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xcaravel_hack_soc_175 la_data_out[47] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_124_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xcaravel_hack_soc_153 la_data_out[24] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xcaravel_hack_soc_164 la_data_out[36] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_124_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xcaravel_hack_soc_186 la_data_out[58] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xcaravel_hack_soc_197 wbs_dat_o[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_3_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_49_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_52_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4830_ _2202_ _0224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_18_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1790 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4761_ soc.rom_encoder_0.request_data_out\[7\] _1481_ _2155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_53_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6500_ _0373_ clknet_leaf_49_wb_clk_i soc.ram_encoder_0.request_data_out\[13\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4692_ soc.spi_video_ram_1.state_sram_clk_counter\[5\] _2104_ _2096_ _2107_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_14_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3712_ _1279_ _1305_ _1309_ _1276_ _1310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_6431_ _0304_ clknet_leaf_78_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[3\]\[17\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3643_ _1222_ _1240_ _1241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_127_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6362_ _0235_ clknet_leaf_132_wb_clk_i soc.spi_video_ram_1.write_fifo.read_pointer\[2\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5313_ soc.ram_encoder_0.request_data_out\[2\] _2545_ _2548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3574_ _1155_ _1157_ _1161_ _1171_ _1172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XFILLER_142_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6293_ _0168_ clknet_leaf_89_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[4\]\[22\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5244_ _1489_ _2495_ _2496_ _0344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_114_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5175_ _2436_ _2442_ _0329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4126_ soc.rom_encoder_0.output_buffer\[4\] _1671_ _1672_ soc.rom_encoder_0.request_address\[3\]
+ _1673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_68_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4057_ _1578_ _1610_ _1613_ _0039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_71_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_52_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4959_ soc.rom_encoder_0.data_out\[14\] soc.rom_encoder_0.request_data_out\[14\]
+ _2287_ _2290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_138_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6629_ soc.cpu.PC.in\[12\] net88 soc.cpu.AReg.data\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_20_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_10_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_16_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_124_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3290_ soc.cpu.ALU.no _0901_ _0902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XTAP_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5931_ _2955_ _0572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_80_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5862_ soc.ram_encoder_0.address\[9\] soc.cpu.AReg.data\[9\] _2902_ _2913_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_90_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5793_ soc.cpu.PC.REG.data\[5\] _2863_ _2864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_4813_ soc.spi_video_ram_1.fifo_in_address\[1\] soc.cpu.AReg.data\[1\] _2018_ _2194_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4744_ _2122_ _2141_ _2142_ _0198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_30_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4675_ soc.spi_video_ram_1.state_sram_clk_counter\[0\] _2094_ _2095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_6414_ _0287_ clknet_leaf_10_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[3\]\[0\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3626_ _1158_ _1159_ _1224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_6345_ _0219_ clknet_leaf_75_wb_clk_i soc.spi_video_ram_1.fifo_in_address\[4\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_3557_ soc.boot_loading_offset\[3\] _1155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_143_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6276_ _0151_ clknet_leaf_124_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[4\]\[5\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_115_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3488_ _1067_ _1083_ _1089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_5227_ _1406_ _2380_ _2482_ _2483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_131_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_88_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5158_ _2400_ _2429_ _0325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_29_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4109_ _1652_ _1645_ _1657_ _0047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_45_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5089_ soc.spi_video_ram_1.write_fifo.fifo_mem\[3\]\[24\] soc.spi_video_ram_1.fifo_in_address\[8\]
+ _2368_ _2375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_16_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_53_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_8_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_15_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4460_ _1961_ _1969_ _1970_ _0085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_3411_ _1010_ _1015_ _1016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4391_ soc.spi_video_ram_1.write_fifo.fifo_mem\[2\]\[22\] soc.spi_video_ram_1.write_fifo.fifo_mem\[3\]\[22\]
+ _1584_ _1914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_131_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3342_ _0853_ _0950_ _0951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_6130_ _0010_ clknet_leaf_8_wb_clk_i net65 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_113_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3273_ _0850_ soc.cpu.ALU.x\[1\] _0885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6061_ soc.spi_video_ram_1.write_fifo.fifo_mem\[2\]\[4\] soc.spi_video_ram_1.fifo_in_data\[4\]
+ _3020_ _3025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_85_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5012_ _2327_ _0281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_38_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5914_ soc.gpio_i_stored\[0\] _2943_ _2861_ _2944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_81_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5845_ _0855_ _2903_ _2904_ _0537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_50_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5776_ _2845_ _2851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_108_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4727_ _2122_ _2128_ _2129_ _0194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_108_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4658_ soc.spi_video_ram_1.write_fifo.fifo_mem\[4\]\[24\] soc.spi_video_ram_1.fifo_in_address\[8\]
+ _2057_ _2084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3609_ soc.video_generator_1.h_count\[3\] soc.video_generator_1.h_count\[4\] _1207_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_66_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4589_ _1933_ _2026_ _2047_ _0137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_6328_ _0203_ clknet_leaf_23_wb_clk_i soc.rom_encoder_0.output_buffer\[15\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6259_ _0134_ clknet_leaf_85_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[7\]\[17\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_103_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_72_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_68_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_79_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3960_ _1529_ _1530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_63_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_50_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3891_ _1190_ _1466_ _1131_ _1469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5630_ _2761_ _0464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_78_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5561_ soc.spi_video_ram_1.fifo_in_data\[12\] soc.spi_video_ram_1.write_fifo.fifo_mem\[5\]\[12\]
+ _2719_ _2721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_117_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5492_ _2436_ _2599_ _0413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4512_ _0009_ _0902_ _2005_ _0102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_144_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4443_ _0688_ _0726_ _0735_ _1958_ _1959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_4374_ soc.spi_video_ram_1.output_buffer\[9\] _1612_ _1899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6113_ _3051_ _3052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_3325_ _0926_ _0934_ _0935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3256_ soc.cpu.AReg.data\[14\] soc.cpu.AReg.data\[13\] _0869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XTAP_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6044_ soc.spi_video_ram_1.fifo_in_address\[10\] soc.spi_video_ram_1.write_fifo.fifo_mem\[1\]\[26\]
+ _2985_ _3015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_67_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3187_ soc.spi_video_ram_1.output_buffer\[18\] _0801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_2309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5828_ soc.cpu.PC.REG.data\[11\] soc.cpu.PC.REG.data\[12\] soc.cpu.PC.REG.data\[13\]
+ _2881_ _2890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_50_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5759_ _0878_ _0902_ _0920_ _0942_ _2835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_10_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_5_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_116_wb_clk_i clknet_4_8_0_wb_clk_i clknet_leaf_116_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_110_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3110_ _0726_ _0728_ _0691_ _0006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4090_ _1497_ _1634_ _1642_ _0043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_95_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_36_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6800_ _0642_ clknet_leaf_108_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[2\]\[13\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_36_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4992_ _2272_ _2312_ _2313_ _0275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_56_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3943_ soc.ram_encoder_0.initializing_step\[0\] _1494_ _1516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6731_ _0573_ clknet_leaf_129_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[0\]\[2\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3874_ _1132_ _1249_ _1455_ _1457_ _1458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
X_6662_ _0504_ clknet_leaf_98_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[6\]\[14\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_118_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5613_ soc.rom_loader.current_address\[1\] _2744_ soc.rom_loader.current_address\[2\]
+ _2750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_20_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6593_ net31 clknet_leaf_24_wb_clk_i soc.rom_encoder_0.data_out\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5544_ soc.spi_video_ram_1.fifo_in_data\[4\] soc.spi_video_ram_1.write_fifo.fifo_mem\[5\]\[4\]
+ _2705_ _2712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_118_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5475_ _1493_ _1490_ _1495_ _2663_ _2664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_144_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4426_ _1592_ _1942_ _1945_ _1702_ _1946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_99_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_101_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4357_ _1761_ _1878_ _1881_ _1882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_101_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3308_ _0916_ _0918_ soc.cpu.ALU.f _0919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4288_ soc.spi_video_ram_1.write_fifo.fifo_mem\[4\]\[10\] soc.spi_video_ram_1.write_fifo.fifo_mem\[5\]\[10\]
+ soc.spi_video_ram_1.write_fifo.fifo_mem\[6\]\[10\] soc.spi_video_ram_1.write_fifo.fifo_mem\[7\]\[10\]
+ _1755_ _1590_ _1817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_104_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3239_ _0849_ _0851_ _0852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_6027_ _3006_ _0617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2117 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2106 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2139 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2128 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xfanout87 net88 net87 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_70_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_2_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_18_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1961 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1950 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1994 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1983 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1972 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3590_ _1130_ _1133_ _1187_ _1188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_115_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5260_ net2 _2505_ _2508_ _2509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_141_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4211_ _1595_ soc.spi_video_ram_1.write_fifo.fifo_mem\[6\]\[5\] _1744_ _1711_ _1745_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_96_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5191_ _2390_ _2454_ _2455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4142_ _1522_ _1681_ _1682_ _0055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_110_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4073_ soc.spi_video_ram_1.write_fifo.fifo_mem\[7\]\[17\] _1628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_110_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_84_wb_clk_i clknet_4_14_0_wb_clk_i clknet_leaf_84_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_110_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xclkbuf_leaf_13_wb_clk_i clknet_4_3_0_wb_clk_i clknet_leaf_13_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_37_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_64_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4975_ _2293_ _2300_ _2301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_52_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3926_ soc.ram_encoder_0.output_bits_left\[4\] _1498_ _1499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_6714_ _0556_ clknet_leaf_8_wb_clk_i soc.boot_loading_offset\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_137_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6645_ _0487_ net90 soc.cpu.ALU.x\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3857_ _1413_ _1443_ _1444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6576_ _0449_ clknet_leaf_105_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[5\]\[24\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3788_ _0759_ _0763_ _1379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_118_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5527_ _2691_ _2700_ _0423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_133_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5458_ _2522_ _2624_ _2625_ _2650_ _2651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_105_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5389_ soc.ram_encoder_0.toggled_sram_sck _1491_ _2595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_99_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4409_ soc.spi_video_ram_1.write_fifo.fifo_mem\[5\]\[20\] _1930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_8_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_129_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xcaravel_hack_soc_121 io_out[26] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xcaravel_hack_soc_110 io_oeb[35] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xcaravel_hack_soc_132 la_data_out[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xcaravel_hack_soc_143 la_data_out[14] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xcaravel_hack_soc_165 la_data_out[37] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_124_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xcaravel_hack_soc_154 la_data_out[25] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xcaravel_hack_soc_176 la_data_out[48] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_123_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xcaravel_hack_soc_198 wbs_dat_o[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xcaravel_hack_soc_187 la_data_out[59] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_105_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_78_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1791 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1780 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4760_ _2122_ _2153_ _2154_ _0202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_61_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4691_ soc.spi_video_ram_1.state_sram_clk_counter\[5\] _2104_ _2106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_3711_ _1306_ _1308_ _1279_ _1309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_6430_ _0303_ clknet_leaf_80_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[3\]\[16\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3642_ _1208_ _1212_ _1213_ _1240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
Xclkbuf_leaf_131_wb_clk_i clknet_4_2_0_wb_clk_i clknet_leaf_131_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_60_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6361_ _0234_ clknet_leaf_132_wb_clk_i soc.spi_video_ram_1.write_fifo.read_pointer\[1\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_143_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5312_ soc.ram_encoder_0.data_out\[2\] _2547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3573_ _1166_ _1169_ _1170_ _1171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
X_6292_ _0167_ clknet_leaf_96_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[4\]\[21\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5243_ soc.ram_encoder_0.input_bits_left\[2\] _2494_ _2496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5174_ _0887_ _2393_ _2441_ _2442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_69_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4125_ _1651_ _1670_ _1672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_60_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_84_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4056_ soc.spi_video_ram_1.output_buffer\[1\] _1612_ _1613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_65_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4958_ _2289_ _0265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_24_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4889_ net6 _2243_ _1955_ _2246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3909_ _1479_ _1483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6628_ soc.cpu.PC.in\[11\] net88 soc.cpu.AReg.data\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_20_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6559_ _0432_ clknet_leaf_120_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[5\]\[7\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_105_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_71_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5930_ soc.spi_video_ram_1.write_fifo.fifo_mem\[0\]\[1\] soc.spi_video_ram_1.fifo_in_data\[1\]
+ _2953_ _2955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_18_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5861_ _2912_ _0545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_61_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5792_ soc.cpu.PC.REG.data\[4\] _2859_ _2863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_4812_ _2193_ _0215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4743_ soc.rom_encoder_0.output_buffer\[10\] _2138_ _2142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_30_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6413_ _0286_ clknet_leaf_44_wb_clk_i net61 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4674_ net69 _2093_ _2094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3625_ _1214_ _1221_ _1222_ _1223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_115_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6344_ _0218_ clknet_leaf_75_wb_clk_i soc.spi_video_ram_1.fifo_in_address\[3\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_3556_ _1147_ _1152_ _1153_ soc.boot_loading_offset\[3\] _1154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_142_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6275_ _0150_ clknet_leaf_124_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[4\]\[4\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_103_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3487_ _1018_ _1019_ _1078_ _1088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5226_ _2480_ _2478_ _2482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_130_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5157_ _0926_ _2392_ _2428_ _2429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_96_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4108_ _1652_ _1656_ _1645_ _1657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_56_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5088_ _2374_ _0310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_29_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4039_ _1584_ _1596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_38_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_53_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_138_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_4_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_133_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_16_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3410_ _0853_ _1014_ _1015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4390_ soc.spi_video_ram_1.write_fifo.fifo_mem\[0\]\[22\] soc.spi_video_ram_1.write_fifo.fifo_mem\[1\]\[22\]
+ _1584_ _1913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_124_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3341_ _0948_ _0949_ _0950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3272_ _0883_ _0884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6060_ _3024_ _0632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5011_ _2326_ soc.rom_encoder_0.request_address\[13\] _2271_ _2327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_23_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5913_ _2942_ _2943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_53_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5844_ soc.ram_encoder_0.address\[0\] _2903_ _2904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_61_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5775_ soc.cpu.PC.REG.data\[0\] soc.cpu.PC.REG.data\[1\] _2850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_108_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4726_ soc.rom_encoder_0.output_buffer\[6\] _1670_ _1672_ soc.rom_encoder_0.request_address\[5\]
+ _2129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4657_ _2083_ _0169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3608_ _1203_ _1205_ _1206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6327_ _0202_ clknet_leaf_23_wb_clk_i soc.rom_encoder_0.output_buffer\[14\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4588_ soc.spi_video_ram_1.fifo_in_address\[4\] _2023_ _2047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_143_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3539_ soc.hack_wait_clocks\[1\] soc.hack_wait_clocks\[0\] _1136_ _0741_ _1137_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_27_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_131_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6258_ _0133_ clknet_leaf_86_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[7\]\[16\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_76_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5209_ _1656_ _2465_ _2469_ _0676_ _0336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_6189_ _0069_ clknet_leaf_110_wb_clk_i soc.spi_video_ram_1.output_buffer\[11\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_29_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_12_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_121_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_44_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3890_ _1190_ _1466_ _1468_ _0018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_43_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5560_ _2720_ _0436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5491_ _2675_ _0412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xclkbuf_leaf_38_wb_clk_i clknet_4_7_0_wb_clk_i clknet_leaf_38_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_89_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4511_ soc.spi_video_ram_1.fifo_in_data\[1\] _2003_ _2005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4442_ _0708_ _0705_ _0732_ soc.spi_video_ram_1.current_state\[4\] _1958_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_99_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_113_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4373_ _0729_ _1877_ _1897_ _1898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_113_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6112_ _2894_ _2919_ _3051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_3324_ _0887_ soc.cpu.AReg.data\[3\] _0928_ _0933_ _0894_ _0934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
XFILLER_86_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3255_ soc.cpu.AReg.data\[0\] _0864_ _0866_ _0868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_58_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6043_ _3014_ _0625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_85_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3186_ soc.spi_video_ram_1.output_buffer\[19\] _0800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_81_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_23_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5827_ _2847_ _2888_ _2889_ _2849_ _0533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_10_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5758_ _0990_ _1091_ _2834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_120_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4709_ soc.spi_video_ram_1.state_sram_clk_counter\[8\] _2116_ soc.spi_video_ram_1.sram_sck_fall_edge
+ soc.spi_video_ram_1.current_state\[4\] _2117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
X_5689_ _1669_ _2779_ _2796_ _0489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_2_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_100_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_60_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4991_ soc.rom_encoder_0.request_address\[7\] _2272_ _2313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_64_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_56_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6730_ _0572_ clknet_leaf_127_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[0\]\[1\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3942_ _1491_ _1496_ _1515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_44_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_3873_ _1268_ _1456_ _1457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6661_ _0503_ clknet_leaf_88_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[6\]\[13\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6592_ net30 clknet_leaf_34_wb_clk_i soc.rom_encoder_0.data_out\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5612_ _2749_ _0458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5543_ _2711_ _0428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_9_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_144_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5474_ _1492_ _2594_ _2663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4425_ _1596_ soc.spi_video_ram_1.write_fifo.fifo_mem\[6\]\[19\] _1944_ _1591_ _1945_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_63_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4356_ _1580_ _1880_ _1881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_87_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3307_ _0917_ _0906_ _0915_ _0918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_140_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4287_ _1814_ _1815_ _1580_ _1816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3238_ _0850_ soc.cpu.ALU.x\[0\] _0851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6026_ soc.spi_video_ram_1.fifo_in_address\[1\] soc.spi_video_ram_1.write_fifo.fifo_mem\[1\]\[17\]
+ _2999_ _3006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2107 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3169_ _0750_ _0783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XTAP_2129 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2118 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout88 soc.cpu.AReg.clk net88 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_136_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1940 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1951 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1995 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1984 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1973 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1962 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_139_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4210_ _1585_ _1743_ _1744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5190_ _1426_ _1420_ _2454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_122_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4141_ soc.ram_encoder_0.output_buffer\[2\] _1509_ _1682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_96_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_68_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4072_ _1601_ soc.spi_video_ram_1.write_fifo.fifo_mem\[4\]\[17\] _1626_ _1627_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_23_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4974_ soc.cpu.PC.REG.data\[3\] _2300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_24_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3925_ soc.ram_encoder_0.output_bits_left\[2\] _1497_ _1498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_leaf_53_wb_clk_i clknet_4_12_0_wb_clk_i clknet_leaf_53_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_51_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6713_ _0555_ clknet_leaf_8_wb_clk_i soc.boot_loading_offset\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6644_ _0486_ net90 soc.cpu.ALU.x\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_20_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3856_ soc.rom_encoder_0.output_buffer\[17\] _1417_ _1442_ soc.rom_encoder_0.request_data_out\[13\]
+ _1443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_20_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3787_ _1378_ net71 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_118_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6575_ _0448_ clknet_leaf_104_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[5\]\[23\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_20_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5526_ _2687_ _2698_ _2700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_132_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5457_ soc.ram_encoder_0.request_data_out\[12\] _2605_ _2650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_106_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4408_ soc.spi_video_ram_1.write_fifo.fifo_mem\[0\]\[20\] soc.spi_video_ram_1.write_fifo.fifo_mem\[1\]\[20\]
+ soc.spi_video_ram_1.write_fifo.fifo_mem\[2\]\[20\] soc.spi_video_ram_1.write_fifo.fifo_mem\[3\]\[20\]
+ _1594_ _1588_ _1929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_120_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5388_ soc.ram_encoder_0.initializing_step\[3\] _2592_ _2593_ _2594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_87_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4339_ _1862_ _1864_ _1865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_86_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6009_ soc.spi_video_ram_1.fifo_in_data\[9\] _2986_ _2997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_55_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_82_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_23_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_10_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xcaravel_hack_soc_100 io_oeb[8] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_6_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xcaravel_hack_soc_111 io_oeb[36] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xcaravel_hack_soc_122 io_out[30] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_137_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xcaravel_hack_soc_155 la_data_out[26] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xcaravel_hack_soc_166 la_data_out[38] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xcaravel_hack_soc_133 la_data_out[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xcaravel_hack_soc_144 la_data_out[15] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xcaravel_hack_soc_177 la_data_out[49] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xcaravel_hack_soc_199 wbs_dat_o[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xcaravel_hack_soc_188 la_data_out[60] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_78_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1792 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1781 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3710_ _1261_ _1307_ _1286_ _1308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4690_ _2104_ _2105_ _0180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3641_ _1223_ _1228_ _1239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_6360_ _0233_ clknet_leaf_132_wb_clk_i soc.spi_video_ram_1.write_fifo.read_pointer\[0\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3572_ _1125_ _1139_ _1128_ _1164_ _1170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_114_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5311_ _2544_ _2542_ _2546_ _0361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_53_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6291_ _0166_ clknet_leaf_119_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[4\]\[20\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_130_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5242_ soc.ram_encoder_0.input_bits_left\[2\] _2494_ _2495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_102_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_100_wb_clk_i clknet_4_10_0_wb_clk_i clknet_leaf_100_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_102_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5173_ _2260_ _2413_ _2414_ _2440_ _2441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_69_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4124_ _1670_ _1671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_60_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput1 io_in[10] net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_57_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4055_ _1611_ _1612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_37_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4957_ soc.rom_encoder_0.data_out\[13\] soc.rom_encoder_0.request_data_out\[13\]
+ _2287_ _2289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4888_ soc.rom_encoder_0.input_buffer\[1\] _2245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3908_ _1478_ _1434_ _1421_ _1482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_137_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6627_ soc.cpu.PC.in\[10\] net88 soc.cpu.AReg.data\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_3839_ soc.rom_encoder_0.current_state\[2\] _1426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_6558_ _0431_ clknet_leaf_81_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[5\]\[6\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_20_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_106_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6489_ _0362_ clknet_leaf_63_wb_clk_i soc.ram_encoder_0.request_data_out\[2\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5509_ soc.hack_clock_0.counter\[4\] _2687_ soc.hack_clock_0.counter\[6\] _2688_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_86_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_2_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5860_ soc.ram_encoder_0.address\[8\] soc.cpu.AReg.data\[8\] _2902_ _2912_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_74_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4811_ soc.spi_video_ram_1.fifo_in_address\[0\] soc.cpu.AReg.data\[0\] _2018_ _2193_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_2290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5791_ _2846_ _2860_ _2862_ _0524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_61_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4742_ soc.rom_encoder_0.request_address\[9\] _1650_ _2125_ soc.rom_encoder_0.output_buffer\[6\]
+ _2140_ _2141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_21_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4673_ soc.spi_video_ram_1.state_counter\[0\] _2091_ _2092_ _2093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6412_ _0285_ clknet_leaf_44_wb_clk_i net60 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3624_ _1212_ _1213_ _1208_ _1222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_115_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6343_ _0217_ clknet_leaf_78_wb_clk_i soc.spi_video_ram_1.fifo_in_address\[2\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_3555_ _1151_ _1149_ _1150_ _1153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_131_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3486_ _1080_ _1084_ _1086_ _1087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_6274_ _0149_ clknet_leaf_123_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[4\]\[3\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5225_ soc.rom_encoder_0.initializing_step\[3\] _2476_ _2481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_84_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5156_ _2252_ _2413_ _2414_ _2427_ _2428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_5_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4107_ _1408_ _1435_ _1656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_56_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5087_ soc.spi_video_ram_1.write_fifo.fifo_mem\[3\]\[23\] soc.spi_video_ram_1.fifo_in_address\[7\]
+ _2368_ _2374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_29_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4038_ _1594_ _1595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_71_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_53_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5989_ _2985_ _2986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_21_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_20_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_4_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_63_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_30_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3340_ _0887_ soc.cpu.AReg.data\[4\] _0894_ _0949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_140_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3271_ _0882_ _0883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5010_ soc.cpu.PC.REG.data\[13\] soc.rom_loader.current_address\[13\] _2292_ _2326_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_94_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5912_ _0744_ _0867_ _2942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_34_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5843_ _2902_ _2903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_34_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_22_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5774_ soc.cpu.PC.REG.data\[0\] _2846_ _2848_ _2849_ _0520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_4725_ soc.rom_encoder_0.output_buffer\[2\] _2125_ _2128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4656_ soc.spi_video_ram_1.write_fifo.fifo_mem\[4\]\[23\] soc.spi_video_ram_1.fifo_in_address\[7\]
+ _2057_ _2083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3607_ _1175_ _1204_ _1205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_4587_ _1943_ _2026_ _2046_ _0136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_6326_ _0201_ clknet_leaf_24_wb_clk_i soc.rom_encoder_0.output_buffer\[13\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3538_ soc.rom_encoder_0.initialized _1136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_107_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3469_ _0884_ _1069_ _1070_ soc.cpu.PC.in\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_6257_ _0132_ clknet_leaf_93_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[7\]\[15\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_88_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5208_ _1419_ _2468_ soc.rom_encoder_0.current_state\[1\] _2469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6188_ _0068_ clknet_leaf_110_wb_clk_i soc.spi_video_ram_1.output_buffer\[12\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_84_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5139_ soc.rom_encoder_0.request_data_out\[4\] _2395_ _2415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_29_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_84_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_8_wb_clk_i clknet_4_1_0_wb_clk_i clknet_leaf_8_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_80_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_138_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_107_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_4_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5490_ _2490_ _2670_ _2671_ _1493_ _0690_ _2675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_4510_ _0009_ _0878_ _2004_ _0101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_8_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4441_ _1957_ _0079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xclkbuf_leaf_78_wb_clk_i clknet_4_14_0_wb_clk_i clknet_leaf_78_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6111_ _3050_ _0657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4372_ _0686_ _1882_ _1896_ _1850_ _1897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_112_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3323_ _0929_ _0868_ _0932_ _0933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3254_ _0855_ _0864_ _0866_ _0867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_86_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_86_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6042_ soc.spi_video_ram_1.fifo_in_address\[9\] soc.spi_video_ram_1.write_fifo.fifo_mem\[1\]\[25\]
+ _2985_ _3014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_67_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3185_ soc.spi_video_ram_1.output_buffer\[17\] _0799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_39_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_96_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5826_ soc.cpu.PC.in\[13\] _2851_ _2889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5757_ _0922_ _1057_ _2833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_22_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4708_ _0682_ _2115_ _2116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_108_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5688_ soc.cpu.ALU.x\[15\] _2777_ _2796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_135_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4639_ _2074_ _0160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_89_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6309_ _0184_ clknet_leaf_137_wb_clk_i soc.spi_video_ram_1.state_sram_clk_counter\[8\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffnq_2
XFILLER_131_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_125_wb_clk_i clknet_4_3_0_wb_clk_i clknet_leaf_125_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_4990_ _2293_ soc.rom_loader.current_address\[7\] _2311_ _2312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_64_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3941_ _1513_ _1514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_56_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6660_ _0502_ clknet_leaf_91_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[6\]\[12\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_17_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3872_ soc.video_generator_1.h_count\[4\] _1131_ _1456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5611_ soc.rom_loader.current_address\[1\] _2744_ _2748_ _2749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_83_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6591_ net28 clknet_leaf_94_wb_clk_i soc.rom_encoder_0.data_out\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5542_ soc.spi_video_ram_1.fifo_in_data\[3\] soc.spi_video_ram_1.write_fifo.fifo_mem\[5\]\[3\]
+ _2705_ _2711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_118_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5473_ _2534_ _2601_ _2662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_8_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4424_ _1756_ _1943_ _1944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_99_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4355_ _1879_ _1880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_101_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3306_ _0852_ _0874_ _0896_ _0899_ _0886_ _0917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_2
XFILLER_58_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4286_ soc.spi_video_ram_1.write_fifo.fifo_mem\[4\]\[28\] soc.spi_video_ram_1.write_fifo.fifo_mem\[5\]\[28\]
+ soc.spi_video_ram_1.write_fifo.fifo_mem\[6\]\[28\] soc.spi_video_ram_1.write_fifo.fifo_mem\[7\]\[28\]
+ _1755_ _1590_ _1815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_101_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_100_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3237_ soc.cpu.ALU.zx _0850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_6025_ _3005_ _0616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2108 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3168_ _0762_ _0768_ _0774_ _0778_ _0781_ _0782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XTAP_2119 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3099_ soc.spi_video_ram_1.state_sram_clk_counter\[7\] soc.spi_video_ram_1.current_state\[4\]
+ _0716_ _0718_ _0719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
Xfanout89 net91 net89 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_5809_ soc.cpu.PC.REG.data\[9\] _2875_ _2876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_50_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6789_ _0631_ clknet_leaf_10_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[2\]\[2\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_13_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_77_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1941 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1952 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1930 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1985 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1974 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1963 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1996 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4140_ soc.ram_encoder_0.request_address\[1\] _1514_ _1681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_68_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4071_ _1596_ _1625_ _1626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_83_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_83_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4973_ _2299_ _0270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_51_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3924_ soc.ram_encoder_0.output_bits_left\[3\] _1497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6712_ _0554_ clknet_leaf_6_wb_clk_i soc.hack_rom_request vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6643_ _0485_ net90 soc.cpu.ALU.x\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_20_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3855_ _1417_ _1437_ _1442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
Xclkbuf_leaf_93_wb_clk_i clknet_4_15_0_wb_clk_i clknet_leaf_93_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_118_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6574_ _0447_ clknet_leaf_89_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[5\]\[22\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3786_ _0807_ _1377_ _1378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_30_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5525_ _2691_ _2698_ _2699_ _0422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
Xclkbuf_leaf_22_wb_clk_i clknet_4_4_0_wb_clk_i clknet_leaf_22_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_5456_ _2615_ _2649_ _0403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4407_ _1686_ _1927_ _1928_ _0074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_132_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5387_ soc.ram_encoder_0.initializing_step\[1\] soc.ram_encoder_0.initializing_step\[0\]
+ _2593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_99_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4338_ _1710_ _1863_ _1579_ _1864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_87_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4269_ soc.spi_video_ram_1.write_fifo.fifo_mem\[1\]\[9\] _1799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_74_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6008_ _1781_ _2988_ _2996_ _0608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_82_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_126_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_7_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xcaravel_hack_soc_123 io_out[31] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xcaravel_hack_soc_112 io_oeb[37] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xcaravel_hack_soc_101 io_oeb[9] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_136_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xcaravel_hack_soc_145 la_data_out[16] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xcaravel_hack_soc_156 la_data_out[28] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xcaravel_hack_soc_134 la_data_out[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_3_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xcaravel_hack_soc_178 la_data_out[50] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xcaravel_hack_soc_189 la_data_out[61] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xcaravel_hack_soc_167 la_data_out[39] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_78_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_78_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1760 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1793 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1782 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1771 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3640_ _1203_ _1205_ _1237_ _1238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_128_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3571_ _1167_ _1168_ _1169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_5310_ soc.ram_encoder_0.request_data_out\[1\] _2545_ _2546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6290_ _0165_ clknet_leaf_87_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[4\]\[19\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_127_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5241_ _0674_ _2493_ _2494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_46_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5172_ soc.rom_encoder_0.request_data_out\[12\] _2394_ _2440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_96_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_96_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4123_ _0674_ _1410_ _1431_ _1670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
Xclkbuf_leaf_140_wb_clk_i clknet_4_2_0_wb_clk_i clknet_leaf_140_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
Xinput2 io_in[11] net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
X_4054_ _0689_ _0705_ _1576_ _1611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_2
XFILLER_28_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_37_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4956_ _2288_ _0264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_40_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4887_ _2240_ _2242_ _2244_ _0239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3907_ _1418_ _1481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_20_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6626_ soc.cpu.PC.in\[9\] net87 soc.cpu.AReg.data\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3838_ soc.rom_encoder_0.initializing_step\[4\] soc.rom_encoder_0.initializing_step\[3\]
+ soc.rom_encoder_0.initializing_step\[2\] soc.rom_encoder_0.initializing_step\[1\]
+ _1425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or4_1
X_6557_ _0430_ clknet_leaf_122_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[5\]\[5\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_118_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5508_ soc.hack_clock_0.counter\[5\] _2687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3769_ _1125_ _1169_ _1336_ _1361_ net74 vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_6488_ _0361_ clknet_leaf_58_wb_clk_i soc.ram_encoder_0.request_data_out\[1\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_126_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5439_ soc.ram_data_out\[7\] _2603_ _2636_ _2637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_106_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_4_6_0_wb_clk_i clknet_0_wb_clk_i clknet_4_6_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_71_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_16_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4810_ soc.spi_video_ram_1.state_sram_clk_counter\[8\] _2116_ _0729_ _0214_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_22_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_33_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5790_ soc.cpu.PC.in\[4\] _2847_ _2861_ _2862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_15_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4741_ soc.rom_encoder_0.request_data_out\[2\] _1481_ _2140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_4672_ _2091_ _1962_ _2092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_135_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6411_ _0284_ clknet_leaf_59_wb_clk_i net59 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3623_ _1215_ _1220_ _1221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6342_ _0216_ clknet_leaf_76_wb_clk_i soc.spi_video_ram_1.fifo_in_address\[1\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_3554_ _1149_ _1150_ _1151_ _1152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_143_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3485_ _1085_ _1086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6273_ _0148_ clknet_leaf_14_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[4\]\[2\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_115_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5224_ soc.rom_encoder_0.initializing_step\[3\] _2480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_97_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5155_ soc.rom_encoder_0.request_data_out\[8\] _2394_ _2427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_57_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4106_ _1415_ _1645_ _1655_ _0046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_57_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5086_ _2373_ _0309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_25_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4037_ _1593_ _1594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_37_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5988_ _2984_ _2985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
X_4939_ _2279_ _0256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_36_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6609_ _0466_ clknet_leaf_29_wb_clk_i soc.rom_loader.current_address\[9\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_125_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_opt_1_0_wb_clk_i clknet_4_0_0_wb_clk_i clknet_opt_1_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_4_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_56_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_15_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3270_ soc.cpu.instruction\[15\] soc.cpu.instruction\[5\] _0882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_87_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5911_ net14 _2941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_59_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5842_ _2901_ _2902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_50_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5773_ _0743_ _2849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_61_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4724_ _2122_ _2126_ _2127_ _0193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_30_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4655_ _2082_ _0168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3606_ _1154_ _1172_ _1166_ _1204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4586_ soc.spi_video_ram_1.fifo_in_address\[3\] _2023_ _2046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6325_ _0200_ clknet_leaf_24_wb_clk_i soc.rom_encoder_0.output_buffer\[12\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3537_ soc.video_generator_1.h_count\[9\] _1134_ _1135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_131_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3468_ _0846_ soc.cpu.ALU.zx soc.cpu.AReg.data\[11\] _0881_ _1070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_6256_ _0131_ clknet_leaf_88_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[7\]\[14\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_97_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3399_ _0979_ _1000_ _0999_ _1004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_69_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5207_ _2389_ _2462_ _2463_ _2468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_6187_ _0067_ clknet_leaf_115_wb_clk_i soc.spi_video_ram_1.output_buffer\[13\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_112_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_111_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5138_ _2391_ _2414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_57_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5069_ _2364_ _0301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_73_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_52_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_75_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_17_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4440_ _1955_ _1956_ _1957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_125_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_113_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6110_ soc.spi_video_ram_1.write_fifo.fifo_mem\[2\]\[28\] soc.spi_video_ram_1.fifo_in_address\[12\]
+ _3019_ _3050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4371_ _0703_ _1888_ _1895_ _1896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_140_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3322_ net80 _0931_ _0867_ soc.gpio_i_stored\[3\] _0868_ _0932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XTAP_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3253_ _0865_ _0866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_79_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6041_ _3013_ _0624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xclkbuf_leaf_47_wb_clk_i clknet_4_6_0_wb_clk_i clknet_leaf_47_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3184_ _0762_ _0795_ _0797_ _0798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_113_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5825_ soc.cpu.PC.REG.data\[13\] _2887_ _2888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_5756_ _0922_ _1038_ _2832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_50_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5687_ _1123_ _2779_ _2795_ _0488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4707_ soc.spi_video_ram_1.state_sram_clk_counter\[2\] soc.spi_video_ram_1.state_sram_clk_counter\[1\]
+ soc.spi_video_ram_1.state_sram_clk_counter\[3\] _2115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4638_ soc.spi_video_ram_1.write_fifo.fifo_mem\[4\]\[14\] soc.spi_video_ram_1.fifo_in_data\[14\]
+ _2069_ _2074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_116_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4569_ _2022_ _2037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_6308_ _0183_ clknet_leaf_137_wb_clk_i soc.spi_video_ram_1.state_sram_clk_counter\[7\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffnq_2
XFILLER_134_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_89_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6239_ _0114_ clknet_leaf_75_wb_clk_i soc.spi_video_ram_1.fifo_in_data\[13\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XTAP_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_41_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3940_ _1493_ _1511_ _1512_ _1513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_91_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3871_ _1190_ _1296_ _1455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_31_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6590_ net27 clknet_4_13_0_wb_clk_i soc.rom_encoder_0.data_out\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5610_ soc.rom_loader.current_address\[1\] _2744_ _2745_ _2748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_13_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5541_ _2710_ _0427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_31_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5472_ _2471_ _2661_ _0407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_144_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4423_ soc.spi_video_ram_1.write_fifo.fifo_mem\[7\]\[19\] _1943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_141_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4354_ soc.spi_video_ram_1.write_fifo.fifo_mem\[4\]\[24\] soc.spi_video_ram_1.write_fifo.fifo_mem\[5\]\[24\]
+ soc.spi_video_ram_1.write_fifo.fifo_mem\[6\]\[24\] soc.spi_video_ram_1.write_fifo.fifo_mem\[7\]\[24\]
+ _1582_ _0001_ _1879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_113_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3305_ _0906_ _0915_ _0916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_98_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6024_ soc.spi_video_ram_1.fifo_in_address\[0\] soc.spi_video_ram_1.write_fifo.fifo_mem\[1\]\[16\]
+ _2999_ _3005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4285_ soc.spi_video_ram_1.write_fifo.fifo_mem\[0\]\[28\] soc.spi_video_ram_1.write_fifo.fifo_mem\[1\]\[28\]
+ soc.spi_video_ram_1.write_fifo.fifo_mem\[2\]\[28\] soc.spi_video_ram_1.write_fifo.fifo_mem\[3\]\[28\]
+ _1755_ _1590_ _1814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_3236_ soc.cpu.ALU.nx _0849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XTAP_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_104_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3167_ _0780_ _0781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_2109 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_54_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3098_ soc.spi_video_ram_1.state_sram_clk_counter\[6\] soc.spi_video_ram_1.state_sram_clk_counter\[5\]
+ soc.spi_video_ram_1.state_sram_clk_counter\[4\] _0717_ _0718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_27_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_82_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_23_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5808_ soc.cpu.PC.REG.data\[8\] _2872_ _2875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_22_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6788_ _0630_ clknet_leaf_128_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[2\]\[1\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_109_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_10_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5739_ _2823_ _0512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_109_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1942 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1920 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1986 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1975 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1964 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1953 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1997 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4070_ soc.spi_video_ram_1.write_fifo.fifo_mem\[5\]\[17\] _1625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_95_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4972_ _2298_ soc.rom_encoder_0.request_address\[2\] _2287_ _2299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_17_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3923_ soc.ram_encoder_0.current_state\[1\] _1488_ _1496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_6711_ _0553_ clknet_leaf_49_wb_clk_i soc.ram_step1_write_request vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6642_ _0484_ net90 soc.cpu.ALU.x\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3854_ _1437_ _1440_ _1441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_20_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_20_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6573_ _0446_ clknet_leaf_95_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[5\]\[21\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_9_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3785_ _1362_ _1368_ _1372_ _1375_ _1376_ _1377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_117_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5524_ soc.hack_clock_0.counter\[4\] _2696_ _2699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_106_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5455_ soc.ram_data_out\[11\] _2604_ _2648_ _2649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xclkbuf_leaf_62_wb_clk_i clknet_4_13_0_wb_clk_i clknet_leaf_62_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_4406_ soc.spi_video_ram_1.output_buffer\[6\] _1611_ _1928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5386_ soc.ram_encoder_0.initializing_step\[4\] soc.ram_encoder_0.initializing_step\[2\]
+ _2592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_113_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4337_ soc.spi_video_ram_1.write_fifo.fifo_mem\[2\]\[13\] soc.spi_video_ram_1.write_fifo.fifo_mem\[3\]\[13\]
+ _1582_ _1863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_101_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4268_ soc.spi_video_ram_1.write_fifo.fifo_mem\[2\]\[9\] soc.spi_video_ram_1.write_fifo.fifo_mem\[3\]\[9\]
+ _1593_ _1798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_74_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3219_ soc.spi_video_ram_1.output_buffer\[4\] _0833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6007_ soc.spi_video_ram_1.fifo_in_data\[8\] _2986_ _2996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4199_ _0800_ _1686_ _1722_ _1733_ _0061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_27_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_126_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_109_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xcaravel_hack_soc_102 io_oeb[14] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xcaravel_hack_soc_113 io_out[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xcaravel_hack_soc_157 la_data_out[29] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xcaravel_hack_soc_146 la_data_out[17] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xcaravel_hack_soc_135 la_data_out[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xcaravel_hack_soc_124 io_out[32] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xcaravel_hack_soc_179 la_data_out[51] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xcaravel_hack_soc_168 la_data_out[40] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_2_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_105_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_3_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_65_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1761 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1750 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1794 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1783 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1772 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_42_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3570_ soc.video_generator_1.v_count\[7\] _1126_ _1127_ _1168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_143_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_143_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5240_ _1501_ _2489_ _2492_ _2493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_142_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5171_ _2436_ _2439_ _0328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_39_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4122_ _1658_ _0881_ _1669_ _0848_ _0048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_68_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4053_ _1581_ _1589_ _1606_ _1609_ _1610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
Xinput3 io_in[12] net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_37_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_101_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4955_ soc.rom_encoder_0.data_out\[12\] soc.rom_encoder_0.request_data_out\[12\]
+ _2287_ _2288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_80_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3906_ soc.rom_encoder_0.output_buffer\[16\] _1440_ _1479_ _1480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_4886_ net5 _2243_ _1955_ _2244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_32_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6625_ soc.cpu.PC.in\[8\] net88 soc.cpu.AReg.data\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3837_ _1411_ _1418_ _1423_ _1424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_118_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6556_ _0429_ clknet_leaf_13_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[5\]\[4\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3768_ soc.video_generator_1.v_count\[8\] soc.video_generator_1.v_count\[1\] _1361_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_5507_ soc.hack_clock_0.counter\[0\] _2686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_69_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6487_ _0360_ clknet_leaf_55_wb_clk_i soc.ram_encoder_0.request_data_out\[0\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3699_ soc.video_generator_1.h_count\[1\] _1216_ _1218_ _1297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5438_ _2512_ _2624_ _2625_ _2635_ _2636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_5369_ _2583_ _0382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_59_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_143_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_81_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4740_ _2122_ _2137_ _2139_ _0197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_14_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4671_ soc.spi_video_ram_1.current_state\[3\] _0703_ soc.spi_video_ram_1.current_state\[0\]
+ soc.spi_video_ram_1.current_state\[2\] _2091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_128_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6410_ _0283_ clknet_leaf_42_wb_clk_i net58 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3622_ _1217_ _1218_ _1219_ _1220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_6341_ _0215_ clknet_leaf_79_wb_clk_i soc.spi_video_ram_1.fifo_in_address\[0\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_127_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3553_ soc.boot_loading_offset\[2\] _1151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_89_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3484_ _1072_ _1075_ _1085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_6272_ _0147_ clknet_leaf_128_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[4\]\[1\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_6_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5223_ _2383_ _2472_ _2477_ _2479_ _0690_ _0340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_116_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5154_ _2400_ _2426_ _0324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_84_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4105_ _1646_ _1648_ _1651_ _1654_ _1655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_29_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5085_ soc.spi_video_ram_1.write_fifo.fifo_mem\[3\]\[22\] soc.spi_video_ram_1.fifo_in_address\[6\]
+ _2368_ _2373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4036_ _1583_ _1593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_38_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_53_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5987_ _0700_ _2703_ _0698_ _2984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_40_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4938_ soc.rom_encoder_0.data_out\[4\] soc.rom_encoder_0.request_data_out\[4\] _2276_
+ _2279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_36_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4869_ _2225_ _2228_ _1403_ _2229_ _2230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_6608_ _0465_ clknet_leaf_30_wb_clk_i soc.rom_loader.current_address\[8\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_20_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6539_ _0412_ clknet_leaf_40_wb_clk_i soc.ram_encoder_0.current_state\[2\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_4_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_29_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_31_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_119_wb_clk_i clknet_4_9_0_wb_clk_i clknet_leaf_119_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_121_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5910_ _0942_ _2936_ _2940_ _0566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_35_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5841_ _2896_ _2899_ _2901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_62_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_22_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5772_ soc.cpu.PC.in\[0\] _2847_ _2848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_50_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_15_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4723_ soc.rom_encoder_0.output_buffer\[5\] _1670_ _1672_ soc.rom_encoder_0.request_address\[4\]
+ _2127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_21_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4654_ soc.spi_video_ram_1.write_fifo.fifo_mem\[4\]\[22\] soc.spi_video_ram_1.fifo_in_address\[6\]
+ _2057_ _2082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4585_ _1618_ _2025_ _2045_ _0135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3605_ _1193_ _1199_ _1203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_6324_ _0199_ clknet_leaf_25_wb_clk_i soc.rom_encoder_0.output_buffer\[11\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3536_ _1130_ _1133_ _1134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_116_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6255_ _0130_ clknet_leaf_88_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[7\]\[13\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_115_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3467_ _0922_ _1060_ _1068_ _1069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
X_5206_ _2436_ _2467_ _0335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_112_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_3398_ _0884_ _1002_ _1003_ soc.cpu.PC.in\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_6186_ _0066_ clknet_leaf_113_wb_clk_i soc.spi_video_ram_1.output_buffer\[14\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_111_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5137_ _2394_ _2413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_29_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5068_ soc.spi_video_ram_1.write_fifo.fifo_mem\[3\]\[14\] soc.spi_video_ram_1.fifo_in_data\[14\]
+ _2357_ _2364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_72_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4019_ _0674_ _0706_ _0188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_16_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_4_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_88_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_76_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4370_ _1710_ _1891_ _1894_ _1579_ _1895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_113_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3321_ soc.cpu.AReg.data\[0\] _0864_ _0930_ _0931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XTAP_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3252_ soc.cpu.AReg.data\[3\] soc.cpu.AReg.data\[2\] soc.cpu.AReg.data\[1\] _0865_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XTAP_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6040_ soc.spi_video_ram_1.fifo_in_address\[8\] soc.spi_video_ram_1.write_fifo.fifo_mem\[1\]\[24\]
+ _2985_ _3013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_26_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_140_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3183_ _0765_ _0796_ _0797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_21_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_87_wb_clk_i clknet_4_9_0_wb_clk_i clknet_leaf_87_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_19_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_16_wb_clk_i clknet_4_6_0_wb_clk_i clknet_leaf_16_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_50_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5824_ soc.cpu.PC.REG.data\[11\] soc.cpu.PC.REG.data\[12\] _2881_ _2887_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_23_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5755_ net84 _2691_ _2831_ _0519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_31_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5686_ soc.cpu.ALU.x\[14\] _2777_ _2795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4706_ _2114_ _0187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_108_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4637_ _2073_ _0159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_144_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4568_ _2036_ _0127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_2_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3519_ _1094_ _1087_ _1100_ _1118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6307_ _0182_ clknet_leaf_137_wb_clk_i soc.spi_video_ram_1.state_sram_clk_counter\[6\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
X_4499_ _1126_ _1995_ soc.video_generator_1.v_count\[7\] _1997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_6238_ _0113_ clknet_leaf_74_wb_clk_i soc.spi_video_ram_1.fifo_in_data\[12\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_58_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6169_ _0049_ clknet_leaf_26_wb_clk_i soc.rom_encoder_0.output_buffer\[4\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_21_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_49_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_49_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3870_ _1432_ _1453_ _1454_ _0676_ _0012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_143_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5540_ soc.spi_video_ram_1.fifo_in_data\[2\] soc.spi_video_ram_1.write_fifo.fifo_mem\[5\]\[2\]
+ _2705_ _2710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_9_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5471_ soc.ram_data_out\[15\] _2604_ _2660_ _2661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_69_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xclkbuf_leaf_134_wb_clk_i clknet_4_2_0_wb_clk_i clknet_leaf_134_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_4422_ _1601_ soc.spi_video_ram_1.write_fifo.fifo_mem\[4\]\[19\] _1941_ _1942_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_144_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4353_ soc.spi_video_ram_1.write_fifo.fifo_mem\[0\]\[24\] soc.spi_video_ram_1.write_fifo.fifo_mem\[1\]\[24\]
+ soc.spi_video_ram_1.write_fifo.fifo_mem\[2\]\[24\] soc.spi_video_ram_1.write_fifo.fifo_mem\[3\]\[24\]
+ _1755_ _1590_ _1878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_87_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3304_ _0853_ _0914_ _0915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4284_ _1353_ _1354_ _1813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_3235_ _0845_ soc.cpu.instruction\[5\] _0848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6023_ _3004_ _0615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_67_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3166_ _0752_ _0779_ _0780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_82_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3097_ soc.spi_video_ram_1.state_sram_clk_counter\[3\] _0711_ soc.spi_video_ram_1.state_sram_clk_counter\[0\]
+ _0717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_1409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_23_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3999_ _1556_ _1560_ _1561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5807_ _2846_ _2873_ _2874_ _2849_ _0528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_6787_ _0629_ clknet_leaf_11_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[2\]\[0\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_109_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5738_ soc.spi_video_ram_1.write_fifo.fifo_mem\[6\]\[22\] soc.spi_video_ram_1.fifo_in_address\[6\]
+ _2798_ _2823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_136_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5669_ _0970_ _2778_ _2786_ _0479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_116_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_2_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_45_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1910 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_54_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1932 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1943 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1921 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1976 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1965 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1954 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1998 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1987 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_127_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_126_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_76_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_64_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4971_ soc.cpu.PC.REG.data\[2\] soc.rom_loader.current_address\[2\] _2293_ _2298_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3922_ _1488_ _1494_ _1495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_6710_ _0552_ clknet_leaf_39_wb_clk_i soc.ram_step2_read_request vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_32_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6641_ _0483_ net90 soc.cpu.ALU.x\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3853_ _1438_ _1439_ _1440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_20_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3784_ _1364_ _1362_ _1376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6572_ _0445_ clknet_leaf_119_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[5\]\[20\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5523_ soc.hack_clock_0.counter\[4\] _2696_ _2698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_30_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5454_ _2520_ _2624_ _2625_ _2647_ _2648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_105_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5385_ _2591_ _0390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_114_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4405_ _1140_ _1921_ _1926_ _1609_ _1927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_87_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4336_ _1756_ soc.spi_video_ram_1.write_fifo.fifo_mem\[0\]\[13\] _1861_ _1862_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_114_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4267_ _1797_ _0065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xclkbuf_leaf_31_wb_clk_i clknet_4_5_0_wb_clk_i clknet_leaf_31_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_3218_ soc.spi_video_ram_1.buffer_index\[4\] _0823_ _0831_ _0832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_28_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4198_ _1581_ _1729_ _1732_ _1720_ _1733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_6006_ _1775_ _2988_ _2995_ _0607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3149_ soc.spi_video_ram_1.buffer_index\[0\] soc.spi_video_ram_1.buffer_index\[1\]
+ _0763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_82_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xcaravel_hack_soc_103 io_oeb[15] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xcaravel_hack_soc_114 io_out[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xcaravel_hack_soc_147 la_data_out[18] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_124_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xcaravel_hack_soc_136 la_data_out[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xcaravel_hack_soc_125 io_out[33] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xcaravel_hack_soc_169 la_data_out[41] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xcaravel_hack_soc_158 la_data_out[30] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_123_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_78_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_19_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1751 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1740 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1784 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1773 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1762 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1795 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_127_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5170_ soc.cpu.ALU.zx _2393_ _2438_ _2439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_110_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4121_ _0990_ _1661_ _1668_ _1669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
XFILLER_69_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4052_ _0710_ _1608_ _1609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_110_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput4 io_in[13] net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_65_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4954_ _2271_ _2287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_3905_ _1419_ _1478_ _1479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4885_ _2241_ _2243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_33_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6624_ soc.cpu.PC.in\[7\] net88 soc.cpu.AReg.data\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3836_ _1416_ _1421_ _1422_ _1403_ _1423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_20_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6555_ _0428_ clknet_leaf_15_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[5\]\[3\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3767_ _1328_ _1189_ _1359_ _1360_ net75 vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
X_5506_ _2681_ _2685_ _0417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_106_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6486_ _0359_ clknet_leaf_49_wb_clk_i soc.ram_encoder_0.request_write vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3698_ soc.video_generator_1.h_count\[3\] soc.video_generator_1.h_count\[2\] _1296_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5437_ soc.ram_encoder_0.request_data_out\[7\] _2606_ _2635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_105_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5368_ soc.ram_encoder_0.address\[6\] soc.ram_encoder_0.request_address\[6\] _2581_
+ _2583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5299_ _2536_ _2537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_59_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4319_ soc.spi_video_ram_1.write_fifo.fifo_mem\[4\]\[26\] soc.spi_video_ram_1.write_fifo.fifo_mem\[5\]\[26\]
+ soc.spi_video_ram_1.write_fifo.fifo_mem\[6\]\[26\] soc.spi_video_ram_1.write_fifo.fifo_mem\[7\]\[26\]
+ _1582_ _1586_ _1846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_101_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4670_ _2090_ _0175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3621_ soc.video_generator_1.h_count\[2\] _1196_ _1219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_30_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6340_ _0214_ clknet_leaf_141_wb_clk_i soc.spi_video_ram_1.sram_sio_oe vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3552_ _1142_ soc.video_generator_1.v_count\[2\] soc.video_generator_1.v_count\[1\]
+ _1143_ _1150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_51_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_142_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3483_ _1067_ _1083_ _1084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6271_ _0146_ clknet_leaf_14_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[4\]\[0\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5222_ _1406_ _2380_ _2478_ _2479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_96_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5153_ _0954_ _2392_ _2425_ _2426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_116_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4104_ _1433_ _1653_ _1654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5084_ _2372_ _0308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_65_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4035_ _1591_ _1592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_80_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_53_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5986_ _2983_ _0599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4937_ _2278_ _0255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_52_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_36_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4868_ soc.rom_encoder_0.request_write _1417_ _2222_ _2229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6607_ _0464_ clknet_leaf_30_wb_clk_i soc.rom_loader.current_address\[7\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3819_ soc.rom_encoder_0.current_state\[0\] _1406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
X_4799_ _2176_ _2184_ _2186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_115_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6538_ _0411_ clknet_leaf_38_wb_clk_i soc.ram_encoder_0.current_state\[1\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_4
XFILLER_107_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6469_ _0342_ clknet_leaf_8_wb_clk_i soc.rom_encoder_0.initializing_step\[4\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_106_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_88_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_62_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5840_ _2897_ _2900_ _0536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_61_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2090 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_99_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5771_ _2845_ _2847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_61_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4722_ soc.rom_encoder_0.output_buffer\[1\] _2125_ _2126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xinput40 la_data_in[4] net40 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_4653_ _2081_ _0167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4584_ soc.spi_video_ram_1.fifo_in_address\[2\] _2023_ _2045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3604_ _1176_ _1186_ _1201_ _1202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_116_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6323_ _0198_ clknet_leaf_23_wb_clk_i soc.rom_encoder_0.output_buffer\[10\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3535_ soc.video_generator_1.h_count\[5\] _1131_ _1132_ _1133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_143_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3466_ _0954_ _1066_ _1067_ _1068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_89_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6254_ _0129_ clknet_leaf_91_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[7\]\[12\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5205_ _1419_ _2466_ _2467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_3397_ _0845_ _0954_ soc.cpu.AReg.data\[7\] _0881_ _1003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_85_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6185_ _0065_ clknet_leaf_135_wb_clk_i soc.spi_video_ram_1.output_buffer\[15\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_97_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5136_ _2400_ _2412_ _0320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5067_ _2363_ _0300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_84_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4018_ _1573_ _1574_ _1575_ _1576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_26_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5969_ soc.spi_video_ram_1.write_fifo.fifo_mem\[0\]\[20\] soc.spi_video_ram_1.fifo_in_address\[4\]
+ _2952_ _2975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_139_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_122_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3320_ soc.cpu.AReg.data\[1\] _0861_ _0930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_113_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3251_ _0856_ _0857_ _0858_ _0859_ _0864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_67_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3182_ _0776_ soc.spi_video_ram_1.output_buffer\[20\] _0772_ soc.spi_video_ram_1.output_buffer\[21\]
+ _0796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_26_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_27_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5823_ _2847_ _2885_ _2886_ _2849_ _0532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_34_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_56_wb_clk_i clknet_4_12_0_wb_clk_i clknet_leaf_56_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_5754_ net84 _0535_ _2831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5685_ _1108_ _2779_ _2794_ _0487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4705_ net69 _2093_ _2096_ _2114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_31_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4636_ soc.spi_video_ram_1.write_fifo.fifo_mem\[4\]\[13\] soc.spi_video_ram_1.fifo_in_data\[13\]
+ _2069_ _2073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_118_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4567_ soc.spi_video_ram_1.fifo_in_data\[10\] soc.spi_video_ram_1.write_fifo.fifo_mem\[7\]\[10\]
+ _2023_ _2036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6306_ _0181_ clknet_leaf_138_wb_clk_i soc.spi_video_ram_1.state_sram_clk_counter\[5\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_144_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3518_ _1096_ _1099_ _1117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4498_ _1126_ _1995_ _1996_ _1984_ _0097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_104_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_3449_ _1026_ _1050_ _1051_ _1052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_6237_ _0112_ clknet_leaf_74_wb_clk_i soc.spi_video_ram_1.fifo_in_data\[11\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_6168_ _0048_ net89 soc.cpu.AReg.data\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_76_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5119_ soc.cpu.DMuxJMP.sel\[0\] _2392_ _2398_ _2399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_58_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_17_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6099_ _3044_ _0651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_45_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_31_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5470_ _2528_ _2606_ _2602_ _2659_ _2660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_9_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4421_ _1585_ _1940_ _1941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_99_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4352_ _1331_ _1877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_98_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3303_ _0907_ _0908_ _0909_ _0913_ soc.cpu.ALU.zy _0914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
Xclkbuf_leaf_103_wb_clk_i clknet_4_10_0_wb_clk_i clknet_leaf_103_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_4283_ _1810_ _1811_ _1812_ _0066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_140_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3234_ soc.cpu.DMuxJMP.sel\[0\] _0847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6022_ soc.spi_video_ram_1.fifo_in_data\[15\] soc.spi_video_ram_1.write_fifo.fifo_mem\[1\]\[15\]
+ _2999_ _3004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_58_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3165_ _0761_ _0779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_39_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3096_ _0715_ _0716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_81_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_70_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3998_ soc.ram_encoder_0.request_data_out\[8\] _1529_ _1557_ _1558_ _1559_ _1560_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_5806_ soc.cpu.PC.in\[8\] _2851_ _2874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6786_ _0628_ clknet_leaf_111_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[1\]\[28\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_10_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5737_ _2822_ _0511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5668_ soc.cpu.ALU.x\[5\] _2784_ _2786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_136_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5599_ _2471_ _2741_ _0454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4619_ soc.spi_video_ram_1.write_fifo.fifo_mem\[4\]\[5\] soc.spi_video_ram_1.fifo_in_data\[5\]
+ _2058_ _2064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_2_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1900 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1933 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1922 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1911 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1977 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1966 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1955 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1944 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1999 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1988 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_139_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_1_wb_clk_i clknet_4_0_0_wb_clk_i clknet_leaf_1_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_126_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4970_ _2297_ _0269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_52_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3921_ soc.ram_encoder_0.initializing_step\[4\] soc.ram_encoder_0.initializing_step\[3\]
+ soc.ram_encoder_0.initializing_step\[2\] soc.ram_encoder_0.initializing_step\[1\]
+ _1494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_6640_ _0482_ net90 soc.cpu.ALU.x\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_60_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3852_ soc.rom_encoder_0.initializing_step\[4\] soc.rom_encoder_0.initializing_step\[3\]
+ soc.rom_encoder_0.initializing_step\[2\] soc.rom_encoder_0.initializing_step\[1\]
+ _1439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_81_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6571_ _0444_ clknet_leaf_87_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[5\]\[19\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5522_ _2691_ _2696_ _2697_ _0421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_3783_ _0809_ _0811_ _0812_ _0815_ _1374_ _1375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_30_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5453_ soc.ram_encoder_0.request_data_out\[11\] _2605_ _2647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_132_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5384_ soc.ram_encoder_0.address\[14\] soc.ram_encoder_0.request_address\[14\] _2581_
+ _2591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4404_ _1922_ _1923_ _1924_ _1925_ _1710_ _1580_ _1926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_99_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4335_ _1593_ _1860_ _1590_ _1861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_59_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4266_ soc.spi_video_ram_1.output_buffer\[15\] _1795_ _1796_ _1797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_67_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3217_ _0808_ _0825_ _0827_ _0811_ _0815_ _0830_ _0831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_6005_ soc.spi_video_ram_1.fifo_in_data\[7\] _2988_ _2995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_39_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4197_ _1605_ _1731_ _1732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_83_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3148_ _0757_ _0760_ _0761_ _0762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XTAP_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3079_ _0697_ _0698_ _0699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_51_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6769_ _0611_ clknet_leaf_95_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[1\]\[11\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_10_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xcaravel_hack_soc_104 io_oeb[20] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_40_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xcaravel_hack_soc_115 io_out[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_137_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xcaravel_hack_soc_126 irq[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xcaravel_hack_soc_148 la_data_out[19] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xcaravel_hack_soc_137 la_data_out[8] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xcaravel_hack_soc_159 la_data_out[31] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_108_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1752 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1730 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_14_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1785 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1763 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1796 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_127_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4120_ _1664_ _1666_ _1667_ _1668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_68_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4051_ soc.spi_video_ram_1.state_sram_clk_counter\[1\] _1607_ _1608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_77_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput5 io_in[16] net5 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_4953_ _2286_ _0263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_91_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3904_ _1407_ soc.rom_encoder_0.current_state\[1\] _1478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_33_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6623_ soc.cpu.PC.in\[6\] net87 soc.cpu.AReg.data\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4884_ _2241_ _2242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_20_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3835_ _1408_ _1419_ _1422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_20_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6554_ _0427_ clknet_leaf_17_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[5\]\[2\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3766_ soc.video_generator_1.h_count\[4\] _1190_ _1131_ _1360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
X_5505_ soc.ram_encoder_0.initializing_step\[4\] _2680_ _2685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_119_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6485_ _0358_ clknet_leaf_46_wb_clk_i soc.ram_encoder_0.input_buffer\[11\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_133_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5436_ _2615_ _2634_ _0398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_10_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3697_ _1277_ _1294_ _1295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_126_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5367_ _2582_ _0381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_142_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5298_ _2490_ _2492_ _2535_ _2536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
X_4318_ soc.spi_video_ram_1.write_fifo.fifo_mem\[0\]\[26\] soc.spi_video_ram_1.write_fifo.fifo_mem\[1\]\[26\]
+ soc.spi_video_ram_1.write_fifo.fifo_mem\[2\]\[26\] soc.spi_video_ram_1.write_fifo.fifo_mem\[3\]\[26\]
+ _1755_ _1587_ _1845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_142_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_102_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4249_ _0802_ _1686_ _1766_ _1780_ _0064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_27_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_82_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_16_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_129_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3620_ soc.video_generator_1.h_count\[1\] _1196_ _1218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_3551_ _1125_ _1128_ _1148_ _1149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_143_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_115_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3482_ _1081_ _1066_ _1082_ _1053_ _1083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_6270_ _0145_ clknet_leaf_117_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[7\]\[28\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_131_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5221_ soc.rom_encoder_0.initializing_step\[2\] soc.rom_encoder_0.initializing_step\[1\]
+ _1438_ _2478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_44_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5152_ _2249_ _2413_ _2414_ _2424_ _2425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_96_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4103_ _1652_ soc.rom_encoder_0.output_bits_left\[3\] _1653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_99_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_96_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5083_ soc.spi_video_ram_1.write_fifo.fifo_mem\[3\]\[21\] soc.spi_video_ram_1.fifo_in_address\[5\]
+ _2368_ _2372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4034_ _1590_ _1591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_64_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5985_ soc.spi_video_ram_1.write_fifo.fifo_mem\[0\]\[28\] soc.spi_video_ram_1.fifo_in_address\[12\]
+ _2952_ _2983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4936_ soc.rom_encoder_0.data_out\[3\] soc.rom_encoder_0.request_data_out\[3\] _2276_
+ _2278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4867_ soc.rom_encoder_0.input_bits_left\[2\] _2226_ _2227_ _2228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_21_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3818_ net81 _1405_ net82 vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6606_ _0463_ clknet_leaf_31_wb_clk_i soc.rom_loader.current_address\[6\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6537_ _0410_ clknet_leaf_38_wb_clk_i soc.ram_encoder_0.current_state\[0\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4798_ _0810_ _2176_ _2184_ _2185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_3749_ soc.spi_video_ram_1.read_value\[2\] soc.spi_video_ram_1.read_value\[3\] _1217_
+ _1347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6468_ _0341_ clknet_leaf_1_wb_clk_i soc.rom_encoder_0.initializing_step\[3\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_5419_ net4 _2488_ _2621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6399_ _0272_ clknet_leaf_27_wb_clk_i soc.rom_encoder_0.request_address\[4\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_121_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_87_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_128_wb_clk_i clknet_4_3_0_wb_clk_i clknet_leaf_128_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_2091 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2080 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5770_ _2845_ _2846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_61_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4721_ _2124_ _2125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_30_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4652_ soc.spi_video_ram_1.write_fifo.fifo_mem\[4\]\[21\] soc.spi_video_ram_1.fifo_in_address\[5\]
+ _2057_ _2081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xinput30 la_data_in[20] net30 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_3603_ _1188_ _1200_ _1201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_116_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4583_ _1628_ _2025_ _2044_ _0134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xinput41 la_data_in[5] net41 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xclkbuf_4_5_0_wb_clk_i clknet_0_wb_clk_i clknet_4_5_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_6322_ _0197_ clknet_leaf_25_wb_clk_i soc.rom_encoder_0.output_buffer\[9\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3534_ soc.video_generator_1.h_count\[7\] _1132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_89_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3465_ _1062_ _1065_ _1067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_6253_ _0128_ clknet_leaf_95_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[7\]\[11\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_103_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5204_ _2230_ _2465_ _2466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_130_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3396_ _0922_ _0992_ _1001_ _1002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
XFILLER_69_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6184_ _0064_ clknet_leaf_113_wb_clk_i soc.spi_video_ram_1.output_buffer\[16\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_96_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5135_ soc.cpu.instruction\[3\] _2392_ _2411_ _2412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5066_ soc.spi_video_ram_1.write_fifo.fifo_mem\[3\]\[13\] soc.spi_video_ram_1.fifo_in_data\[13\]
+ _2357_ _2363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4017_ soc.spi_video_ram_1.state_sram_clk_counter\[1\] _0685_ _1575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_65_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5968_ _2974_ _0590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4919_ soc.rom_encoder_0.input_buffer\[11\] _2266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_138_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5899_ soc.hack_wait_clocks\[1\] _2934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_20_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_99_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3250_ net77 _0855_ _0860_ _0862_ _0863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XTAP_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3181_ _0775_ _0794_ _0795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_78_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5822_ soc.cpu.PC.in\[12\] _2851_ _2886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_22_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5753_ _2830_ _0535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_72_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4704_ net69 _2093_ _2111_ _0186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_5684_ soc.cpu.ALU.x\[13\] _2784_ _2794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_30_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4635_ _2072_ _0158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xclkbuf_leaf_96_wb_clk_i clknet_4_11_0_wb_clk_i clknet_leaf_96_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_116_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_25_wb_clk_i clknet_4_5_0_wb_clk_i clknet_leaf_25_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_4566_ _2035_ _0126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_143_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3517_ _1105_ _1104_ _1115_ _1116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_6305_ _0180_ clknet_leaf_138_wb_clk_i soc.spi_video_ram_1.state_sram_clk_counter\[4\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
X_4497_ _1126_ _1995_ _1996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_131_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3448_ _1029_ _1032_ _1051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6236_ _0111_ clknet_leaf_78_wb_clk_i soc.spi_video_ram_1.fifo_in_data\[10\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_134_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3379_ _0974_ _0978_ _0986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6167_ _0047_ clknet_leaf_4_wb_clk_i soc.rom_encoder_0.output_bits_left\[2\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5118_ _2393_ _2396_ _2397_ _2398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_69_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6098_ soc.spi_video_ram_1.write_fifo.fifo_mem\[2\]\[22\] soc.spi_video_ram_1.fifo_in_address\[6\]
+ _3019_ _3044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_85_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5049_ soc.spi_video_ram_1.write_fifo.fifo_mem\[3\]\[5\] soc.spi_video_ram_1.fifo_in_data\[5\]
+ _2217_ _2354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_80_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_25_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_88_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_20_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_129_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4420_ soc.spi_video_ram_1.write_fifo.fifo_mem\[5\]\[19\] _1940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_8_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4351_ _1811_ _1875_ _1876_ _0070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_141_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3302_ _0868_ _0910_ _0911_ _0912_ _0913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_4_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4282_ soc.spi_video_ram_1.output_buffer\[14\] _1612_ _1812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_101_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3233_ _0845_ _0846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
X_6021_ _1883_ _2988_ _3003_ _0614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_67_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_143_wb_clk_i clknet_opt_1_0_wb_clk_i clknet_leaf_143_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_3164_ _0775_ _0777_ _0778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_95_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_67_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3095_ soc.spi_video_ram_1.state_sram_clk_counter\[8\] _0681_ _0715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_27_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3997_ soc.ram_encoder_0.initializing_step\[0\] _1494_ _1515_ _1559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_5805_ soc.cpu.PC.REG.data\[8\] _2872_ _2873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_50_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6785_ _0627_ clknet_leaf_98_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[1\]\[27\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_22_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5736_ soc.spi_video_ram_1.write_fifo.fifo_mem\[6\]\[21\] soc.spi_video_ram_1.fifo_in_address\[5\]
+ _2798_ _2822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5667_ _0958_ _2778_ _2785_ _0478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_89_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4618_ _2063_ _0150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_117_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5598_ soc.rom_loader.rom_request _2740_ _2268_ _2741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_89_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4549_ soc.spi_video_ram_1.fifo_in_data\[1\] _2026_ _2027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_1_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6219_ _0094_ clknet_leaf_131_wb_clk_i soc.video_generator_1.v_count\[3\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_38_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1901 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1934 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1923 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1967 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1956 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1945 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1989 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1978 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_16_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_64_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3920_ soc.ram_encoder_0.current_state\[2\] _1493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_32_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3851_ soc.rom_encoder_0.initializing_step\[0\] _1438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_20_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6570_ _0443_ clknet_leaf_83_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[5\]\[18\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3782_ _0771_ _1373_ _1374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5521_ soc.hack_clock_0.counter\[3\] _2694_ _2697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_74_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5452_ _2615_ _2646_ _0402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5383_ _2590_ _0389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_99_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4403_ soc.spi_video_ram_1.write_fifo.fifo_mem\[6\]\[21\] soc.spi_video_ram_1.write_fifo.fifo_mem\[7\]\[21\]
+ _1724_ _1925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_99_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4334_ soc.spi_video_ram_1.write_fifo.fifo_mem\[1\]\[13\] _1860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_59_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6004_ _2994_ _0606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4265_ _0689_ _0705_ _1576_ _1796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_86_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4196_ _1730_ _1731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3216_ _0757_ _0828_ _0829_ _0830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_82_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3147_ _0750_ soc.spi_video_ram_1.buffer_index\[1\] _0759_ _0761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_27_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3078_ soc.spi_video_ram_1.write_fifo.write_pointer\[0\] _0698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_36_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_40_wb_clk_i clknet_4_7_0_wb_clk_i clknet_leaf_40_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_6768_ _0610_ clknet_leaf_85_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[1\]\[10\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_7_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6699_ _0541_ clknet_leaf_77_wb_clk_i soc.ram_encoder_0.address\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5719_ _2813_ _0502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xcaravel_hack_soc_105 io_oeb[21] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xcaravel_hack_soc_138 la_data_out[9] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_136_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xcaravel_hack_soc_116 io_out[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xcaravel_hack_soc_127 irq[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xcaravel_hack_soc_149 la_data_out[20] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_105_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_77_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_85_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1742 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1720 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1731 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1775 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1764 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1753 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1797 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1786 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_139_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_127_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_122_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4050_ soc.spi_video_ram_1.state_sram_clk_counter\[8\] soc.spi_video_ram_1.state_sram_clk_counter\[0\]
+ _0684_ _1607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
Xinput6 io_in[17] net6 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_110_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_52_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4952_ soc.rom_encoder_0.data_out\[11\] soc.rom_encoder_0.request_data_out\[11\]
+ _2276_ _2286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_51_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4883_ _1403_ _2223_ _2241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_60_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3903_ soc.rom_encoder_0.initializing_step\[4\] soc.rom_encoder_0.initializing_step\[3\]
+ _1476_ _1477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_6622_ soc.cpu.PC.in\[5\] net87 soc.cpu.AReg.data\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_3834_ soc.rom_encoder_0.current_state\[2\] _1420_ _1421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_60_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6553_ _0426_ clknet_leaf_122_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[5\]\[1\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3765_ soc.video_generator_1.h_count\[4\] _1190_ _1131_ _1359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_5504_ _2684_ _0416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_118_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6484_ _0357_ clknet_leaf_59_wb_clk_i soc.ram_encoder_0.input_buffer\[10\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3696_ _1265_ _1285_ _1293_ _1261_ _1294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_106_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5435_ soc.ram_data_out\[6\] _2603_ _2633_ _2634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_142_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_114_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5366_ soc.ram_encoder_0.address\[5\] soc.ram_encoder_0.request_address\[5\] _2581_
+ _2582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5297_ _1512_ _2533_ _2534_ _2535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_87_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_59_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4317_ _1702_ _1840_ _1843_ _1844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_102_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4248_ _1773_ _1779_ _1780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_142_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4179_ soc.spi_video_ram_1.write_fifo.fifo_mem\[0\]\[2\] soc.spi_video_ram_1.write_fifo.fifo_mem\[1\]\[2\]
+ soc.spi_video_ram_1.write_fifo.fifo_mem\[2\]\[2\] soc.spi_video_ram_1.write_fifo.fifo_mem\[3\]\[2\]
+ _1594_ _1588_ _1716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_71_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_23_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_109_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_133_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_3550_ soc.video_generator_1.v_count\[2\] soc.video_generator_1.v_count\[1\] _1148_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_115_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3481_ _1046_ _1077_ _1082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5220_ soc.rom_encoder_0.initializing_step\[2\] _2476_ _2477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_143_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5151_ soc.rom_encoder_0.request_data_out\[7\] _2395_ _2424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_37_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4102_ soc.rom_encoder_0.output_bits_left\[2\] _1652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5082_ _2371_ _0307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_96_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4033_ _0001_ _1590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_38_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5984_ _2982_ _0598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4935_ _2277_ _0254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_123_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4866_ soc.rom_encoder_0.input_bits_left\[4\] _2227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_20_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3817_ soc.ram_encoder_0.toggled_sram_sck _1405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6605_ _0462_ clknet_leaf_31_wb_clk_i soc.rom_loader.current_address\[5\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4797_ soc.spi_video_ram_1.current_state\[3\] _0764_ _2184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6536_ _0409_ clknet_leaf_40_wb_clk_i soc.ram_encoder_0.sram_sio_oe vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3748_ _1326_ _1188_ _1346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_106_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6467_ _0340_ clknet_leaf_3_wb_clk_i soc.rom_encoder_0.initializing_step\[2\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_3679_ _1264_ _1273_ _1275_ _1239_ _1276_ _1277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_5418_ soc.ram_encoder_0.request_data_out\[3\] _2606_ _2620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_106_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6398_ _0271_ clknet_leaf_27_wb_clk_i soc.rom_encoder_0.request_address\[3\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_121_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5349_ soc.ram_encoder_0.data_out\[14\] _2572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_82_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_43_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_29_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_15_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_120_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2070 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2092 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2081 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4720_ _1412_ _1420_ _1440_ _2123_ _2124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_4651_ _2080_ _0166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput20 la_data_in[11] net20 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput31 la_data_in[21] net31 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_3602_ _1193_ _1199_ _1200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xinput42 la_data_in[6] net42 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_4582_ soc.spi_video_ram_1.fifo_in_address\[1\] _2023_ _2044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_115_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6321_ _0196_ clknet_leaf_25_wb_clk_i soc.rom_encoder_0.output_buffer\[8\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3533_ soc.video_generator_1.h_count\[6\] _1131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_131_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3464_ _1062_ _1065_ _1066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_66_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6252_ _0127_ clknet_leaf_85_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[7\]\[10\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5203_ _2389_ _2462_ _2463_ _2464_ _2465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
X_6183_ _0063_ clknet_leaf_113_wb_clk_i soc.spi_video_ram_1.output_buffer\[17\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_112_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3395_ _0954_ _0999_ _1000_ _1001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5134_ _2393_ _2409_ _2410_ _2411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_85_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5065_ _2362_ _0299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_38_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4016_ soc.spi_video_ram_1.current_state\[4\] _0725_ _0685_ _1574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_25_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5967_ soc.spi_video_ram_1.write_fifo.fifo_mem\[0\]\[19\] soc.spi_video_ram_1.fifo_in_address\[3\]
+ _2964_ _2974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4918_ _2264_ _2243_ _2265_ _0249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_40_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5898_ _2931_ _2933_ _0741_ _0561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_21_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4849_ _0694_ _2213_ _1955_ _2215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_119_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_119_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6519_ _0392_ clknet_leaf_47_wb_clk_i soc.ram_data_out\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_107_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_76_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_7_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3180_ _0776_ soc.spi_video_ram_1.output_buffer\[22\] _0772_ soc.spi_video_ram_1.output_buffer\[23\]
+ _0794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_67_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5821_ soc.cpu.PC.REG.data\[12\] _2884_ _2885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_5752_ _0689_ _2690_ _2830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_50_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4703_ _2093_ _2111_ _0185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5683_ _1092_ _2779_ _2793_ _0486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_30_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4634_ soc.spi_video_ram_1.write_fifo.fifo_mem\[4\]\[12\] soc.spi_video_ram_1.fifo_in_data\[12\]
+ _2069_ _2072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4565_ soc.spi_video_ram_1.fifo_in_data\[9\] soc.spi_video_ram_1.write_fifo.fifo_mem\[7\]\[9\]
+ _2023_ _2035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_144_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_128_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3516_ _1111_ _1114_ _1115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_6304_ _0179_ clknet_leaf_136_wb_clk_i soc.spi_video_ram_1.state_sram_clk_counter\[3\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_103_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4496_ _1984_ _1994_ _1995_ _0096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
Xclkbuf_leaf_65_wb_clk_i clknet_4_12_0_wb_clk_i clknet_leaf_65_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_3447_ _1029_ _1032_ _1050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6235_ _0110_ clknet_leaf_80_wb_clk_i soc.spi_video_ram_1.fifo_in_data\[9\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_3378_ _0979_ _0984_ _0985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_6166_ _0046_ clknet_leaf_4_wb_clk_i soc.rom_encoder_0.output_bits_left\[3\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5117_ net5 _2223_ _2397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6097_ _3043_ _0650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_57_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5048_ _2353_ _0291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_84_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_122_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_88_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_57_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_90_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_32_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_31_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_83_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4350_ soc.spi_video_ram_1.output_buffer\[10\] _1612_ _1876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3301_ soc.cpu.AReg.data\[0\] net39 _0864_ _0866_ _0912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or4_1
XFILLER_140_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4281_ _1575_ _1578_ _1811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_3232_ soc.cpu.instruction\[15\] _0845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_6020_ soc.spi_video_ram_1.fifo_in_data\[14\] _2986_ _3003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_121_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_100_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3163_ _0776_ soc.spi_video_ram_1.output_buffer\[4\] _0772_ soc.spi_video_ram_1.output_buffer\[5\]
+ _0777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_94_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3094_ _0711_ _0713_ _0714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_54_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5804_ _2310_ _2869_ _2872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xclkbuf_leaf_112_wb_clk_i clknet_4_8_0_wb_clk_i clknet_leaf_112_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_23_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3996_ soc.ram_encoder_0.request_write _1558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_22_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6784_ _0626_ clknet_leaf_100_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[1\]\[26\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_31_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5735_ _2821_ _0510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_136_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5666_ soc.cpu.ALU.x\[4\] _2784_ _2785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_30_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4617_ soc.spi_video_ram_1.write_fifo.fifo_mem\[4\]\[4\] soc.spi_video_ram_1.fifo_in_data\[4\]
+ _2058_ _2063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_135_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5597_ soc.rom_loader.wait_fall_clk soc.rom_loader.writing _2738_ _2739_ _2740_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_144_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4548_ _2022_ _2026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_144_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4479_ _1127_ _1167_ _1983_ _0675_ _1984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_4
XFILLER_131_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6218_ _0093_ clknet_leaf_130_wb_clk_i soc.video_generator_1.v_count\[2\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_98_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6149_ _0029_ clknet_leaf_62_wb_clk_i soc.ram_encoder_0.output_buffer\[10\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_86_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1924 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1913 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1902 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_54_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1968 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1957 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1946 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1979 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_139_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_6_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_122_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_76_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3850_ _1427_ _1422_ _1437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_60_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3781_ _0808_ _0814_ _0816_ _0760_ _1373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_13_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5520_ soc.hack_clock_0.counter\[3\] _2694_ _2696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_8_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5451_ soc.ram_data_out\[10\] _2604_ _2645_ _2646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_67_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5382_ soc.ram_encoder_0.address\[13\] soc.ram_encoder_0.request_address\[13\] _2581_
+ _2590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4402_ soc.spi_video_ram_1.write_fifo.fifo_mem\[4\]\[21\] soc.spi_video_ram_1.write_fifo.fifo_mem\[5\]\[21\]
+ _1724_ _1924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_141_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4333_ _1761_ _1855_ _1858_ _1859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_114_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4264_ _1693_ _1695_ _1794_ _1607_ _1795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_6003_ soc.spi_video_ram_1.fifo_in_data\[6\] soc.spi_video_ram_1.write_fifo.fifo_mem\[1\]\[6\]
+ _2986_ _2994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3215_ _0783_ soc.spi_video_ram_1.output_buffer\[21\] _0829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4195_ soc.spi_video_ram_1.write_fifo.fifo_mem\[4\]\[4\] soc.spi_video_ram_1.write_fifo.fifo_mem\[5\]\[4\]
+ soc.spi_video_ram_1.write_fifo.fifo_mem\[6\]\[4\] soc.spi_video_ram_1.write_fifo.fifo_mem\[7\]\[4\]
+ _1593_ _1587_ _1730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_95_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3146_ _0758_ _0759_ _0760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_67_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3077_ soc.spi_video_ram_1.write_fifo.read_pointer\[0\] _0697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_27_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_39_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6767_ _0609_ clknet_leaf_121_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[1\]\[9\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3979_ soc.ram_encoder_0.output_buffer\[12\] _1527_ _1545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5718_ soc.spi_video_ram_1.write_fifo.fifo_mem\[6\]\[12\] soc.spi_video_ram_1.fifo_in_data\[12\]
+ _2810_ _2813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_50_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6698_ _0540_ clknet_leaf_70_wb_clk_i soc.ram_encoder_0.address\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xcaravel_hack_soc_106 io_oeb[27] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_5649_ soc.rom_loader.current_address\[14\] _2773_ _2774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
Xclkbuf_leaf_80_wb_clk_i clknet_4_14_0_wb_clk_i clknet_leaf_80_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
Xcaravel_hack_soc_139 la_data_out[10] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xcaravel_hack_soc_128 irq[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xcaravel_hack_soc_117 io_out[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_104_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_105_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1743 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1721 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1732 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1710 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1776 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1765 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1798 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1787 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_5_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput7 io_in[18] net7 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_64_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_49_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4951_ _2285_ _0262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_36_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4882_ soc.rom_encoder_0.input_buffer\[0\] _2240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3902_ soc.rom_encoder_0.initializing_step\[1\] _1438_ soc.rom_encoder_0.initializing_step\[2\]
+ _1476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6621_ soc.cpu.PC.in\[4\] net87 soc.cpu.AReg.data\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3833_ soc.rom_encoder_0.current_state\[1\] _1419_ _1420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_33_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_20_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6552_ _0425_ clknet_leaf_13_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[5\]\[0\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_9_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3764_ soc.spi_video_ram_1.sram_sio_oe net57 vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_5503_ _2680_ _2683_ _2684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_6483_ _0356_ clknet_leaf_59_wb_clk_i soc.ram_encoder_0.input_buffer\[9\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3695_ _1217_ _1292_ _1276_ _1293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5434_ _2510_ _2624_ _2625_ _2632_ _2633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_114_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5365_ _2537_ _2581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_87_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5296_ _1493_ _1503_ _2534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_102_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4316_ _1761_ _1842_ _1843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_101_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4247_ _1607_ _1778_ _1779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4178_ soc.spi_video_ram_1.output_buffer\[21\] _1715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_83_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3129_ soc.cpu.instruction\[15\] soc.cpu.instruction\[3\] _0744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_82_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6819_ _0661_ clknet_leaf_54_wb_clk_i soc.ram_encoder_0.data_out\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_51_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_27_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_14_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3480_ _1042_ _1045_ _1081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_108_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5150_ _2400_ _2423_ _0323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_111_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4101_ _1650_ _1651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_57_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5081_ soc.spi_video_ram_1.write_fifo.fifo_mem\[3\]\[20\] soc.spi_video_ram_1.fifo_in_address\[4\]
+ _2368_ _2371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4032_ soc.spi_video_ram_1.write_fifo.fifo_mem\[0\]\[16\] soc.spi_video_ram_1.write_fifo.fifo_mem\[1\]\[16\]
+ soc.spi_video_ram_1.write_fifo.fifo_mem\[2\]\[16\] soc.spi_video_ram_1.write_fifo.fifo_mem\[3\]\[16\]
+ _1585_ _1588_ _1589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_110_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5983_ soc.spi_video_ram_1.write_fifo.fifo_mem\[0\]\[27\] soc.spi_video_ram_1.fifo_in_address\[11\]
+ _2952_ _2982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_37_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4934_ soc.rom_encoder_0.data_out\[2\] soc.rom_encoder_0.request_data_out\[2\] _2276_
+ _2277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_40_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_19_wb_clk_i clknet_4_4_0_wb_clk_i clknet_leaf_19_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_4865_ soc.rom_encoder_0.input_bits_left\[3\] _2226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6604_ _0461_ clknet_leaf_32_wb_clk_i soc.rom_loader.current_address\[4\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3816_ net62 _1404_ net63 vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4796_ _0764_ _2177_ _2182_ _2183_ _0209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_6535_ _0408_ clknet_leaf_39_wb_clk_i net81 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_20_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3747_ _1196_ _1249_ _1345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_118_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6466_ _0339_ clknet_leaf_7_wb_clk_i soc.rom_encoder_0.initializing_step\[1\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_3678_ _1230_ _1232_ _1276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_5417_ _2615_ _2619_ _0394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6397_ _0270_ clknet_leaf_27_wb_clk_i soc.rom_encoder_0.request_address\[2\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_133_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5348_ _2570_ _2538_ _2571_ _0373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_130_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5279_ _2520_ _2504_ _2521_ _0354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_102_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_52_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_12_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_59_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_19_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2060 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2093 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2082 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2071 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4650_ soc.spi_video_ram_1.write_fifo.fifo_mem\[4\]\[20\] soc.spi_video_ram_1.fifo_in_address\[4\]
+ _2057_ _2080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xinput21 la_data_in[12] net21 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput10 io_in[23] net10 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_3601_ _1195_ _1198_ _1199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
Xinput32 la_data_in[22] net32 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_6320_ _0195_ clknet_leaf_26_wb_clk_i soc.rom_encoder_0.output_buffer\[7\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xinput43 la_data_in[7] net43 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_4581_ _1602_ _2025_ _2043_ _0133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_116_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_137_wb_clk_i clknet_4_2_0_wb_clk_i clknet_leaf_137_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_3532_ soc.video_generator_1.h_count\[8\] _1130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_3463_ _0926_ _1064_ _1065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_6251_ _0126_ clknet_leaf_81_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[7\]\[9\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_6_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5202_ _1439_ _1428_ _2464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6182_ _0062_ clknet_leaf_114_wb_clk_i soc.spi_video_ram_1.output_buffer\[18\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5133_ net8 _2223_ _2410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3394_ _0994_ _0998_ _1000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_111_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5064_ soc.spi_video_ram_1.write_fifo.fifo_mem\[3\]\[12\] soc.spi_video_ram_1.fifo_in_data\[12\]
+ _2357_ _2362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4015_ soc.spi_video_ram_1.current_state\[3\] soc.spi_video_ram_1.current_state\[0\]
+ _1573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_38_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5966_ _2973_ _0589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_52_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4917_ soc.rom_encoder_0.input_buffer\[6\] _2241_ _2250_ _2265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5897_ soc.hack_wait_clocks\[1\] _2932_ _2933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_34_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4848_ _2213_ _2214_ _0230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_32_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4779_ soc.rom_encoder_0.output_buffer\[14\] _1436_ _2169_ _1441_ _2170_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_119_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6518_ _0391_ clknet_leaf_36_wb_clk_i soc.ram_encoder_0.initialized vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_10_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6449_ _0322_ clknet_leaf_16_wb_clk_i soc.cpu.instruction\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_103_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_34_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5820_ soc.cpu.PC.REG.data\[11\] _2881_ _2884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_35_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_22_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5751_ _2829_ _0518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4702_ _2111_ _2113_ _0184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5682_ soc.cpu.ALU.x\[12\] _2784_ _2793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_30_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4633_ _2071_ _0157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4564_ _1790_ _2025_ _2034_ _0125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_144_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_104_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3515_ _0926_ _1113_ _1114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_6303_ _0178_ clknet_leaf_136_wb_clk_i soc.spi_video_ram_1.state_sram_clk_counter\[2\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_89_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6234_ _0109_ clknet_leaf_80_wb_clk_i soc.spi_video_ram_1.fifo_in_data\[8\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_4495_ _1127_ _1993_ _1995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_3446_ _1005_ _1008_ _1048_ _1049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3377_ _0945_ _0981_ _0983_ _0984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_69_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6165_ _0045_ clknet_leaf_4_wb_clk_i soc.rom_encoder_0.output_bits_left\[4\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5116_ soc.rom_encoder_0.request_data_out\[0\] _2395_ _2396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6096_ soc.spi_video_ram_1.write_fifo.fifo_mem\[2\]\[21\] soc.spi_video_ram_1.fifo_in_address\[5\]
+ _3019_ _3043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5047_ soc.spi_video_ram_1.write_fifo.fifo_mem\[3\]\[4\] soc.spi_video_ram_1.fifo_in_data\[4\]
+ _2217_ _2353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xclkbuf_leaf_34_wb_clk_i clknet_4_7_0_wb_clk_i clknet_leaf_34_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_26_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5949_ soc.spi_video_ram_1.write_fifo.fifo_mem\[0\]\[10\] soc.spi_video_ram_1.fifo_in_data\[10\]
+ _2964_ _2965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_13_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_134_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_75_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_31_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_118_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3300_ soc.gpio_i_stored\[2\] soc.cpu.AReg.data\[0\] _0860_ _0865_ _0911_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_113_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4280_ _0729_ _1356_ _1809_ _1608_ _1810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_113_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3231_ _0844_ net70 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3162_ _0750_ _0776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_67_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_39_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3093_ soc.spi_video_ram_1.state_sram_clk_counter\[3\] _0682_ _0712_ _0713_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_35_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_63_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5803_ _2846_ _2870_ _2871_ _2849_ _0527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_90_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3995_ _1493_ soc.ram_encoder_0.current_state\[1\] _1502_ _1557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_50_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6783_ _0625_ clknet_leaf_106_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[1\]\[25\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_22_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5734_ soc.spi_video_ram_1.write_fifo.fifo_mem\[6\]\[20\] soc.spi_video_ram_1.fifo_in_address\[4\]
+ _2798_ _2821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5665_ _2777_ _2784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_30_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4616_ _2062_ _0149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5596_ soc.rom_encoder_0.write_enable net45 _2739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4547_ _2022_ _2025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_143_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_104_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4478_ soc.video_generator_1.v_count\[2\] _1981_ _1982_ _1983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_132_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3429_ _1029_ _1032_ _1033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_6217_ _0092_ clknet_leaf_131_wb_clk_i soc.video_generator_1.v_count\[1\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_6148_ _0028_ clknet_leaf_63_wb_clk_i soc.ram_encoder_0.output_buffer\[9\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_85_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_73_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6079_ _3034_ _0641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_46_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1925 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1914 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1903 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1958 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1936 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1947 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1969 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_70_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_5_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_1_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_92_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3780_ _0815_ _0839_ _1369_ _1371_ _1372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_5450_ _2518_ _2624_ _2625_ _2644_ _2645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_4401_ soc.spi_video_ram_1.write_fifo.fifo_mem\[2\]\[21\] soc.spi_video_ram_1.write_fifo.fifo_mem\[3\]\[21\]
+ _1724_ _1923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_132_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5381_ _2589_ _0388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_99_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4332_ _1580_ _1857_ _1858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4263_ _1761_ _1783_ _1786_ _1789_ _1793_ _1794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_101_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3214_ soc.spi_video_ram_1.output_buffer\[20\] _0828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6002_ _1734_ _2988_ _2993_ _0605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4194_ soc.spi_video_ram_1.write_fifo.fifo_mem\[0\]\[4\] soc.spi_video_ram_1.write_fifo.fifo_mem\[1\]\[4\]
+ soc.spi_video_ram_1.write_fifo.fifo_mem\[2\]\[4\] soc.spi_video_ram_1.write_fifo.fifo_mem\[3\]\[4\]
+ _1585_ _1711_ _1729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_94_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3145_ soc.spi_video_ram_1.buffer_index\[2\] _0759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_28_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3076_ soc.spi_video_ram_1.write_fifo.read_pointer\[0\] _0693_ _0695_ _0696_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_51_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3978_ soc.ram_encoder_0.output_buffer\[8\] _1520_ _1530_ soc.ram_encoder_0.request_data_out\[4\]
+ _1543_ _1544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_51_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_11_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6766_ _0608_ clknet_leaf_120_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[1\]\[8\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5717_ _2812_ _0501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_108_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6697_ _0539_ clknet_leaf_53_wb_clk_i soc.ram_encoder_0.address\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xcaravel_hack_soc_129 la_data_out[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xcaravel_hack_soc_107 io_oeb[28] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_5648_ soc.rom_loader.current_address\[13\] _2771_ _2773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xcaravel_hack_soc_118 io_out[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_40_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5579_ soc.spi_video_ram_1.fifo_in_address\[5\] soc.spi_video_ram_1.write_fifo.fifo_mem\[5\]\[21\]
+ _2719_ _2730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_2_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_131_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1700 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1722 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1733 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1711 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1766 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1755 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1744 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1799 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1788 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_111_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_39_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_1_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput8 io_in[19] net8 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_76_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4950_ soc.rom_encoder_0.data_out\[10\] soc.rom_encoder_0.request_data_out\[10\]
+ _2276_ _2285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4881_ _2236_ _2239_ _0238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_33_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_3901_ _1460_ _1475_ _0022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6620_ soc.cpu.PC.in\[3\] net87 soc.cpu.AReg.data\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_60_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3832_ _1406_ _1419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_6551_ _0424_ clknet_leaf_38_wb_clk_i soc.hack_clock_0.counter\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5502_ _2681_ _2682_ _2683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3763_ soc.rom_encoder_0.sram_sio_oe net53 vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_6482_ _0355_ clknet_leaf_44_wb_clk_i soc.ram_encoder_0.input_buffer\[8\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3694_ _1286_ _1289_ _1291_ _1292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5433_ soc.ram_encoder_0.request_data_out\[6\] _2606_ _2632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_133_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5364_ _2580_ _0380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4315_ _1841_ _1842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5295_ _2530_ _2532_ _2533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_87_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4246_ _1711_ _1774_ _1777_ _1702_ _1778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_95_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4177_ _0820_ _1686_ _1697_ _1714_ _0058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_83_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3128_ soc.hack_wait_clocks\[1\] soc.hack_wait_clocks\[0\] _0741_ _0742_ _0743_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__or4_1
XFILLER_83_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3059_ _0677_ _0678_ _0679_ _0680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_23_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6818_ _0660_ clknet_leaf_54_wb_clk_i soc.ram_encoder_0.data_out\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_11_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6749_ _0591_ clknet_leaf_118_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[0\]\[20\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_109_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4100_ _1406_ _1478_ _1417_ _1650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
X_5080_ _2370_ _0306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_111_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4031_ _1587_ _1588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_77_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5982_ _2981_ _0597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_80_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4933_ _2271_ _2276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_18_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4864_ _1426_ _2224_ _2225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_32_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_59_wb_clk_i clknet_4_7_0_wb_clk_i clknet_leaf_59_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_6603_ _0460_ clknet_leaf_28_wb_clk_i soc.rom_loader.current_address\[3\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3815_ _1403_ _1404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4795_ _0758_ _2178_ _2183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6534_ _0407_ clknet_leaf_47_wb_clk_i soc.ram_data_out\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3746_ _1318_ _1325_ _1341_ _1343_ _1344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_107_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6465_ _0338_ clknet_leaf_8_wb_clk_i soc.rom_encoder_0.initializing_step\[0\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5416_ soc.ram_data_out\[2\] _2603_ _2618_ _2619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3677_ _1241_ _1274_ _1275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6396_ _0269_ clknet_leaf_27_wb_clk_i soc.rom_encoder_0.request_address\[1\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5347_ soc.ram_encoder_0.request_data_out\[13\] _2566_ _2571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_82_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5278_ soc.ram_encoder_0.input_buffer\[3\] _2505_ _2508_ _2521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_102_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4229_ _1711_ _1754_ _1760_ _1761_ _1762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_75_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2061 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2050 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2094 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2083 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2072 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput11 io_in[24] net11 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_128_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4580_ soc.spi_video_ram_1.fifo_in_address\[0\] _2026_ _2043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xinput22 la_data_in[13] net22 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_3600_ soc.video_generator_1.h_count\[5\] _1197_ _1198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_30_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xinput33 la_data_in[23] net33 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_7_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput44 la_data_in[8] net44 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_3531_ _1125_ _1128_ _1129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_143_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3462_ _1011_ _1063_ _1064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6250_ _0125_ clknet_leaf_121_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[7\]\[8\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3393_ _0994_ _0998_ _0999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5201_ _1406_ _1409_ _2385_ _2463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_6181_ _0061_ clknet_leaf_134_wb_clk_i soc.spi_video_ram_1.output_buffer\[19\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_42_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5132_ soc.rom_encoder_0.request_data_out\[3\] _2395_ _2409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_leaf_106_wb_clk_i clknet_4_10_0_wb_clk_i clknet_leaf_106_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_29_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5063_ _2361_ _0298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4014_ _1522_ _1571_ _1572_ _0038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_65_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_37_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5965_ soc.spi_video_ram_1.write_fifo.fifo_mem\[0\]\[18\] soc.spi_video_ram_1.fifo_in_address\[2\]
+ _2964_ _2973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_34_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4916_ soc.rom_encoder_0.input_buffer\[10\] _2264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5896_ soc.hack_wait_clocks\[0\] _2929_ _2932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4847_ _0698_ _2212_ _1955_ _2214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_119_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4778_ _1413_ _2168_ _2169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6517_ _0390_ clknet_leaf_60_wb_clk_i soc.ram_encoder_0.request_address\[14\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3729_ soc.video_generator_1.h_count\[3\] _1196_ _1220_ _1327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_134_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6448_ _0321_ clknet_leaf_16_wb_clk_i soc.cpu.instruction\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6379_ _0252_ clknet_leaf_21_wb_clk_i soc.rom_encoder_0.request_data_out\[0\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_102_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_102_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_90_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_4_wb_clk_i clknet_4_1_0_wb_clk_i clknet_leaf_4_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_4_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_66_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5750_ soc.spi_video_ram_1.write_fifo.fifo_mem\[6\]\[28\] soc.spi_video_ram_1.fifo_in_address\[12\]
+ _2798_ _2829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5681_ _1069_ _2779_ _2792_ _0485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4701_ soc.spi_video_ram_1.state_sram_clk_counter\[8\] _2112_ _2113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_15_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4632_ soc.spi_video_ram_1.write_fifo.fifo_mem\[4\]\[11\] soc.spi_video_ram_1.fifo_in_data\[11\]
+ _2069_ _2071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_31_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_129_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4563_ soc.spi_video_ram_1.fifo_in_data\[8\] _2026_ _2034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_116_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3514_ _1011_ _1112_ _1113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6302_ _0177_ clknet_leaf_136_wb_clk_i soc.spi_video_ram_1.state_sram_clk_counter\[1\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffnq_2
X_4494_ _1127_ _1993_ _1994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3445_ _1020_ _1034_ _1048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_89_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6233_ _0108_ clknet_leaf_52_wb_clk_i soc.spi_video_ram_1.fifo_in_data\[7\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_6164_ _0044_ clknet_leaf_44_wb_clk_i soc.ram_encoder_0.output_bits_left\[2\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_112_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3376_ _0967_ _0982_ _0983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5115_ _2394_ _2395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_58_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6095_ _3042_ _0649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5046_ _2352_ _0290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_72_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_41_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_74_wb_clk_i clknet_4_15_0_wb_clk_i clknet_leaf_74_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_5948_ _2951_ _2964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_5879_ _1209_ _2739_ _2921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_119_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_88_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_4_4_0_wb_clk_i clknet_0_wb_clk_i clknet_4_4_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_56_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_8_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_8_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_33_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3230_ _0806_ _0807_ _0843_ _0720_ _0844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_140_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3161_ _0751_ _0764_ _0775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_39_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3092_ soc.spi_video_ram_1.state_sram_clk_counter\[8\] soc.spi_video_ram_1.state_sram_clk_counter\[1\]
+ soc.spi_video_ram_1.state_sram_clk_counter\[0\] _0712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_82_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5802_ soc.cpu.PC.in\[7\] _2851_ _2871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_23_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3994_ soc.ram_encoder_0.output_buffer\[12\] _1555_ _1556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6782_ _0624_ clknet_leaf_107_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[1\]\[24\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5733_ _2820_ _0509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5664_ _0942_ _2778_ _2783_ _0477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4615_ soc.spi_video_ram_1.write_fifo.fifo_mem\[4\]\[3\] soc.spi_video_ram_1.fifo_in_data\[3\]
+ _2058_ _2062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5595_ soc.rom_encoder_0.initialized _2268_ _2738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_144_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4546_ _2024_ _0117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_116_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_121_wb_clk_i clknet_4_9_0_wb_clk_i clknet_leaf_121_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_143_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_89_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4477_ _1162_ soc.video_generator_1.v_count\[1\] _1139_ _1982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_104_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3428_ _0853_ _1031_ _1032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_6216_ _0091_ clknet_leaf_9_wb_clk_i soc.video_generator_1.v_count\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6147_ _0027_ clknet_leaf_62_wb_clk_i soc.ram_encoder_0.output_buffer\[8\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3359_ _0962_ _0966_ _0967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_58_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6078_ soc.spi_video_ram_1.write_fifo.fifo_mem\[2\]\[12\] soc.spi_video_ram_1.fifo_in_data\[12\]
+ _3031_ _3034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5029_ _2333_ _2342_ _0283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_38_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1904 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1959 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1948 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1926 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4400_ soc.spi_video_ram_1.write_fifo.fifo_mem\[0\]\[21\] soc.spi_video_ram_1.write_fifo.fifo_mem\[1\]\[21\]
+ _1724_ _1922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_126_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5380_ soc.ram_encoder_0.address\[12\] soc.ram_encoder_0.request_address\[12\] _2581_
+ _2589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4331_ _1856_ _1857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4262_ _1580_ _1792_ _1793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3213_ _0757_ _0801_ _0826_ _0827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6001_ soc.spi_video_ram_1.fifo_in_data\[5\] _2988_ _2993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_79_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4193_ _0828_ _1686_ _1722_ _1728_ _0060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_83_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3144_ soc.spi_video_ram_1.buffer_index\[1\] _0758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_94_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3075_ soc.spi_video_ram_1.write_fifo.read_pointer\[1\] _0694_ _0695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_23_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3977_ soc.ram_encoder_0.request_address\[11\] _1513_ _1543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_11_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6765_ _0607_ clknet_leaf_127_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[1\]\[7\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5716_ soc.spi_video_ram_1.write_fifo.fifo_mem\[6\]\[11\] soc.spi_video_ram_1.fifo_in_data\[11\]
+ _2810_ _2812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6696_ _0538_ clknet_leaf_70_wb_clk_i soc.ram_encoder_0.address\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xcaravel_hack_soc_108 io_oeb[29] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xcaravel_hack_soc_119 io_out[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_5647_ soc.rom_loader.current_address\[13\] _2771_ _2772_ _0470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_3_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5578_ _1930_ _2708_ _2729_ _0445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_116_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4529_ _2003_ _1039_ _2014_ _0110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_144_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1723 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1712 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1701 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1767 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1756 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1745 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1789 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1778 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_10_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_139_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_110_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xinput9 io_in[22] net9 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_76_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_17_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4880_ soc.rom_encoder_0.input_bits_left\[4\] _2237_ _2239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_32_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3900_ soc.video_generator_1.h_count\[9\] _1473_ _1475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_3831_ _1413_ _1417_ _1418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_32_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3762_ soc.ram_encoder_0.sram_sio_oe net49 vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_6550_ _0423_ clknet_leaf_36_wb_clk_i soc.hack_clock_0.counter\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_60_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5501_ soc.ram_encoder_0.initializing_step\[2\] _2678_ soc.ram_encoder_0.initializing_step\[3\]
+ _2682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_72_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_118_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6481_ _0354_ clknet_leaf_46_wb_clk_i soc.ram_encoder_0.input_buffer\[7\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_9_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3693_ _1288_ _1290_ _1269_ _1291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5432_ _2615_ _2631_ _0397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_69_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_127_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5363_ soc.ram_encoder_0.address\[4\] soc.ram_encoder_0.request_address\[4\] _2566_
+ _2580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_126_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4314_ soc.spi_video_ram_1.write_fifo.fifo_mem\[4\]\[12\] soc.spi_video_ram_1.write_fifo.fifo_mem\[5\]\[12\]
+ soc.spi_video_ram_1.write_fifo.fifo_mem\[6\]\[12\] soc.spi_video_ram_1.write_fifo.fifo_mem\[7\]\[12\]
+ _1583_ _1586_ _1841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_114_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5294_ soc.ram_step2_read_request soc.ram_step1_write_request _2531_ _2532_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_101_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4245_ _1596_ _1775_ _1776_ _1591_ _1777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_132_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4176_ _0685_ _1704_ _1713_ _1714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_83_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3127_ soc.ram_encoder_0.initialized soc.rom_encoder_0.initialized soc.spi_video_ram_1.initialized
+ _0742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_71_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3058_ soc.spi_video_ram_1.state_counter\[1\] soc.spi_video_ram_1.state_counter\[0\]
+ soc.spi_video_ram_1.state_counter\[3\] soc.spi_video_ram_1.state_counter\[2\] _0679_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_51_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6817_ _0659_ clknet_leaf_56_wb_clk_i soc.ram_encoder_0.data_out\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_23_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_109_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6748_ _0590_ clknet_leaf_89_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[0\]\[19\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6679_ _0521_ net84 soc.cpu.PC.REG.data\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_118_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_120_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_101_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_127_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4030_ _1586_ _1587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_64_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5981_ soc.spi_video_ram_1.write_fifo.fifo_mem\[0\]\[26\] soc.spi_video_ram_1.fifo_in_address\[10\]
+ _2952_ _2981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_80_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4932_ _2275_ _0253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_64_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_33_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_33_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6602_ _0459_ clknet_leaf_28_wb_clk_i soc.rom_loader.current_address\[2\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_60_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4863_ soc.rom_encoder_0.current_state\[1\] _1406_ _2224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_33_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3814_ soc.rom_encoder_0.toggled_sram_sck _1403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_4794_ _2178_ _2179_ _2182_ _0208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_21_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6533_ _0406_ clknet_leaf_57_wb_clk_i soc.ram_data_out\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3745_ _1342_ _1251_ _1254_ _1343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_20_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6464_ _0337_ clknet_leaf_5_wb_clk_i soc.rom_encoder_0.current_state\[2\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_133_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5415_ _2604_ _2616_ _2617_ _2618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_3676_ _1261_ _1262_ _1274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xclkbuf_leaf_99_wb_clk_i clknet_4_10_0_wb_clk_i clknet_leaf_99_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
Xclkbuf_leaf_28_wb_clk_i clknet_4_5_0_wb_clk_i clknet_leaf_28_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_6395_ _0268_ clknet_leaf_27_wb_clk_i soc.rom_encoder_0.request_address\[0\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_115_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_102_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5346_ soc.ram_encoder_0.data_out\[13\] _2570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5277_ soc.ram_encoder_0.input_buffer\[7\] _2520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_102_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4228_ _1579_ _1761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_29_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4159_ _1685_ _1686_ _1691_ _1697_ _0057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_56_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2040 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2051 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_34_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2095 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2084 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2073 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2062 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xinput12 io_in[25] net12 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput34 la_data_in[24] net34 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput45 la_data_in[9] net45 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput23 la_data_in[14] net23 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_3530_ soc.video_generator_1.v_count\[8\] soc.video_generator_1.v_count\[7\] _1126_
+ _1127_ _1128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_128_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3461_ _0907_ soc.cpu.AReg.data\[11\] _1012_ soc.ram_data_out\[11\] _1063_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_97_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3392_ _0853_ _0997_ _0998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_5200_ _1412_ _1417_ _2459_ _2462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_6180_ _0060_ clknet_leaf_134_wb_clk_i soc.spi_video_ram_1.output_buffer\[20\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_112_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5131_ _2400_ _2408_ _0319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_35_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5062_ soc.spi_video_ram_1.write_fifo.fifo_mem\[3\]\[11\] soc.spi_video_ram_1.fifo_in_data\[11\]
+ _2357_ _2361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4013_ soc.ram_encoder_0.output_buffer\[19\] _1509_ _1572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_111_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_42_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_42_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5964_ _2972_ _0588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_52_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4915_ _2262_ _2242_ _2263_ _0248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_61_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5895_ soc.hack_wait_clocks\[0\] _2929_ _2931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4846_ _0698_ _2212_ _2213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_138_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6516_ _0389_ clknet_leaf_64_wb_clk_i soc.ram_encoder_0.request_address\[13\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4777_ soc.rom_encoder_0.output_buffer\[14\] _1417_ _1442_ soc.rom_encoder_0.request_data_out\[10\]
+ _2168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_20_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3728_ _1193_ _1195_ _1326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6447_ _0320_ clknet_leaf_19_wb_clk_i soc.cpu.instruction\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3659_ _1142_ _1126_ _1257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6378_ _0251_ clknet_leaf_22_wb_clk_i soc.rom_encoder_0.request_write vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5329_ _2557_ _2542_ _2558_ _0367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_103_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5680_ soc.cpu.ALU.x\[11\] _2784_ _2792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4700_ soc.spi_video_ram_1.state_sram_clk_counter\[7\] _2108_ _2112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4631_ _2070_ _0156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_30_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4562_ _1770_ _2025_ _2033_ _0124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_144_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3513_ _0907_ soc.cpu.AReg.data\[14\] _1012_ soc.ram_data_out\[14\] _1112_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6301_ _0176_ clknet_leaf_137_wb_clk_i soc.spi_video_ram_1.state_sram_clk_counter\[0\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffnq_2
X_4493_ _1984_ _1992_ _1993_ _0095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_144_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3444_ _1046_ _1047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6232_ _0107_ clknet_leaf_80_wb_clk_i soc.spi_video_ram_1.fifo_in_data\[6\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_6163_ _0043_ clknet_leaf_42_wb_clk_i soc.ram_encoder_0.output_bits_left\[3\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_112_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3375_ _0947_ _0951_ _0962_ _0966_ _0982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5114_ _2225_ _2394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6094_ soc.spi_video_ram_1.write_fifo.fifo_mem\[2\]\[20\] soc.spi_video_ram_1.fifo_in_address\[4\]
+ _3019_ _3042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5045_ soc.spi_video_ram_1.write_fifo.fifo_mem\[3\]\[3\] soc.spi_video_ram_1.fifo_in_data\[3\]
+ _2217_ _2352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_84_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_72_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5947_ _2963_ _0580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_34_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5878_ _2293_ net45 soc.boot_loading_offset\[0\] _2920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xclkbuf_leaf_43_wb_clk_i clknet_4_7_0_wb_clk_i clknet_leaf_43_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_4829_ soc.spi_video_ram_1.fifo_in_address\[9\] soc.cpu.AReg.data\[9\] _0748_ _2202_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_21_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_17_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3160_ _0765_ _0773_ _0762_ _0774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_79_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3091_ soc.spi_video_ram_1.state_sram_clk_counter\[2\] _0711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_95_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_35_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5801_ soc.cpu.PC.REG.data\[7\] _2869_ _2870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_63_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6781_ _0623_ clknet_leaf_104_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[1\]\[23\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3993_ _1515_ _1518_ _1555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_5732_ soc.spi_video_ram_1.write_fifo.fifo_mem\[6\]\[19\] soc.spi_video_ram_1.fifo_in_address\[3\]
+ _2810_ _2820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5663_ soc.cpu.ALU.x\[3\] _2779_ _2783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_31_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4614_ _2061_ _0148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5594_ _2737_ _0453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_116_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4545_ soc.spi_video_ram_1.fifo_in_data\[0\] soc.spi_video_ram_1.write_fifo.fifo_mem\[7\]\[0\]
+ _2023_ _2024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_143_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4476_ _1125_ soc.video_generator_1.v_count\[8\] soc.video_generator_1.v_count\[7\]
+ _1126_ _1981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_131_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3427_ _1011_ _1030_ _1031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6215_ _0090_ clknet_leaf_143_wb_clk_i soc.spi_video_ram_1.state_counter\[10\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6146_ _0026_ clknet_leaf_67_wb_clk_i soc.ram_encoder_0.output_buffer\[7\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_98_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3358_ _0926_ _0965_ _0966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3289_ _0898_ _0900_ _0901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_6077_ _3033_ _0640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_39_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5028_ _0690_ _2341_ _2342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_85_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1905 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1938 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1949 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1927 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_142_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_21_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_135_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_95_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_103_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_118_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4330_ soc.spi_video_ram_1.write_fifo.fifo_mem\[4\]\[25\] soc.spi_video_ram_1.write_fifo.fifo_mem\[5\]\[25\]
+ soc.spi_video_ram_1.write_fifo.fifo_mem\[6\]\[25\] soc.spi_video_ram_1.write_fifo.fifo_mem\[7\]\[25\]
+ _1582_ _0001_ _1856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_5_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4261_ _1756_ soc.spi_video_ram_1.write_fifo.fifo_mem\[6\]\[8\] _1791_ _1710_ _1792_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_140_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3212_ _0783_ soc.spi_video_ram_1.output_buffer\[19\] _0826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6000_ _2992_ _0604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_79_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4192_ _1581_ _1723_ _1727_ _1720_ _1728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_95_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3143_ _0750_ _0757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_67_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_54_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3074_ soc.spi_video_ram_1.write_fifo.write_pointer\[1\] _0694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_36_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_36_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3976_ _1510_ _1541_ _1542_ _0030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6764_ _0606_ clknet_leaf_14_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[1\]\[6\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_11_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6695_ _0537_ clknet_leaf_53_wb_clk_i soc.ram_encoder_0.address\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5715_ _2811_ _0500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5646_ _2089_ soc.rom_loader.was_loading _2771_ soc.rom_loader.current_address\[13\]
+ _2772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
Xcaravel_hack_soc_109 io_oeb[34] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_117_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5577_ soc.spi_video_ram_1.fifo_in_address\[4\] _2705_ _2729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4528_ soc.spi_video_ram_1.fifo_in_data\[9\] _2007_ _2014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4459_ soc.spi_video_ram_1.state_counter\[5\] _1967_ _1970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_120_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6129_ _1669_ _2896_ _3051_ _2574_ _0673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XTAP_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_86_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1724 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1713 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1702 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_26_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1746 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1735 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1779 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1768 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_76_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_18_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3830_ _1416_ _1417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
X_3761_ _1129_ _1135_ _1358_ net76 vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_32_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5500_ _1488_ _2595_ _0675_ _2681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6480_ _0353_ clknet_leaf_58_wb_clk_i soc.ram_encoder_0.input_buffer\[6\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3692_ _1286_ _1280_ _1290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5431_ soc.ram_data_out\[5\] _2603_ _2630_ _2631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_65_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5362_ _2579_ _0379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_142_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4313_ soc.spi_video_ram_1.write_fifo.fifo_mem\[0\]\[12\] soc.spi_video_ram_1.write_fifo.fifo_mem\[1\]\[12\]
+ soc.spi_video_ram_1.write_fifo.fifo_mem\[2\]\[12\] soc.spi_video_ram_1.write_fifo.fifo_mem\[3\]\[12\]
+ _1724_ _1587_ _1840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_5293_ _0743_ _2531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_141_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4244_ _1756_ soc.spi_video_ram_1.write_fifo.fifo_mem\[0\]\[7\] _1776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4175_ _1592_ _1707_ _1712_ _1605_ _1713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_83_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3126_ soc.rom_encoder_0.write_enable net18 net13 net37 _0741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or4_1
XTAP_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3057_ soc.spi_video_ram_1.state_counter\[5\] soc.spi_video_ram_1.state_counter\[4\]
+ soc.spi_video_ram_1.state_counter\[7\] soc.spi_video_ram_1.state_counter\[6\] _0678_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_42_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6816_ _0658_ clknet_leaf_55_wb_clk_i soc.ram_encoder_0.data_out\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_51_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6747_ _0589_ clknet_leaf_79_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[0\]\[18\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3959_ _1501_ _1511_ _1529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_129_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6678_ _0520_ net84 soc.cpu.PC.REG.data\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_13_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5629_ soc.rom_loader.current_address\[7\] _2759_ _2760_ _2761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_117_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_15_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_30_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_127_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_123_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5980_ _2980_ _0596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_24_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4931_ soc.rom_encoder_0.data_out\[1\] soc.rom_encoder_0.request_data_out\[1\] _2272_
+ _2275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_75_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4862_ _1407_ _1422_ _2223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_6601_ _0458_ clknet_leaf_28_wb_clk_i soc.rom_loader.current_address\[1\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3813_ _1402_ net73 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_33_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4793_ _0689_ _0705_ _2181_ _2182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
X_6532_ _0405_ clknet_leaf_47_wb_clk_i soc.ram_data_out\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3744_ _1247_ _1248_ _1342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_21_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_119_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6463_ _0336_ clknet_leaf_5_wb_clk_i soc.rom_encoder_0.current_state\[1\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_3675_ _1265_ _1267_ _1271_ _1272_ _1273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_127_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5414_ net3 _2488_ _2617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_106_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6394_ _0267_ clknet_leaf_7_wb_clk_i soc.rom_encoder_0.request_data_out\[15\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_114_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5345_ _2568_ _2538_ _2569_ _0372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_99_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5276_ _2518_ _2504_ _2519_ _0353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_114_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4227_ _1591_ _1759_ _1760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_96_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4158_ _1692_ _1578_ _1696_ _1697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_4089_ _1514_ _1634_ _1641_ _1642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_3109_ _0727_ soc.spi_video_ram_1.current_state\[2\] _0728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_28_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_70_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_106_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_121_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_143_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2041 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2052 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2030 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2085 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2074 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2063 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2096 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_122_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xinput13 io_in[26] net13 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput24 la_data_in[15] net24 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput35 la_data_in[25] net35 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_109_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3460_ _0923_ _1061_ _1062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_131_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3391_ _0995_ _0996_ _0997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_111_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5130_ soc.cpu.DMuxJMP.sel\[2\] _2392_ _2407_ _2408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_69_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5061_ _2360_ _0297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_2_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4012_ soc.ram_encoder_0.output_buffer\[15\] _1555_ _1530_ soc.ram_encoder_0.request_data_out\[11\]
+ _1559_ _1571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_42_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5963_ soc.spi_video_ram_1.write_fifo.fifo_mem\[0\]\[17\] soc.spi_video_ram_1.fifo_in_address\[1\]
+ _2964_ _2972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_52_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4914_ soc.rom_encoder_0.input_buffer\[5\] _2241_ _2250_ _2263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_52_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5894_ _2861_ _2929_ _2930_ _0560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_80_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_115_wb_clk_i clknet_4_8_0_wb_clk_i clknet_leaf_115_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_4845_ _1949_ _0740_ _2211_ _2212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4776_ _1671_ _2166_ _2167_ _0205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_21_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6515_ _0388_ clknet_leaf_64_wb_clk_i soc.ram_encoder_0.request_address\[12\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3727_ _1236_ _1324_ _1325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6446_ _0319_ clknet_leaf_16_wb_clk_i soc.cpu.DMuxJMP.sel\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3658_ _1252_ _1254_ _1255_ _1256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_121_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6377_ _0250_ clknet_leaf_18_wb_clk_i soc.rom_encoder_0.input_buffer\[11\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3589_ _1130_ soc.video_generator_1.h_count\[9\] _1133_ _1187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_115_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5328_ soc.ram_encoder_0.request_data_out\[7\] _2545_ _2558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_76_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5259_ _0675_ _2508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_103_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_12_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_11_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4630_ soc.spi_video_ram_1.write_fifo.fifo_mem\[4\]\[10\] soc.spi_video_ram_1.fifo_in_data\[10\]
+ _2069_ _2070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6300_ _0175_ clknet_leaf_22_wb_clk_i soc.rom_loader.was_loading vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4561_ soc.spi_video_ram_1.fifo_in_data\[7\] _2026_ _2033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_128_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3512_ _0923_ _1110_ _1111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_7_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4492_ _1167_ _1991_ _1993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_3443_ _1042_ _1045_ _1046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_6231_ _0106_ clknet_leaf_52_wb_clk_i soc.spi_video_ram_1.fifo_in_data\[5\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_6162_ _0042_ clknet_leaf_42_wb_clk_i soc.ram_encoder_0.output_bits_left\[4\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_103_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3374_ _0980_ _0968_ _0967_ _0981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_5113_ _2391_ _2393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_69_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_58_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6093_ _3041_ _0648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5044_ _2351_ _0289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_81_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5946_ soc.spi_video_ram_1.write_fifo.fifo_mem\[0\]\[9\] soc.spi_video_ram_1.fifo_in_data\[9\]
+ _2953_ _2963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5877_ _2738_ _2919_ _0554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_138_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4828_ _2201_ _0223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_21_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4759_ soc.rom_encoder_0.output_buffer\[14\] _2138_ _2154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_88_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_122_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6429_ _0302_ clknet_leaf_73_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[3\]\[15\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_leaf_83_wb_clk_i clknet_4_9_0_wb_clk_i clknet_leaf_83_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
Xclkbuf_leaf_12_wb_clk_i clknet_4_3_0_wb_clk_i clknet_leaf_12_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_88_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_31_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3090_ _0703_ _0710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_94_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3992_ _1522_ _1553_ _1554_ _0034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5800_ soc.cpu.PC.REG.data\[5\] soc.cpu.PC.REG.data\[6\] _2863_ _2869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_63_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6780_ _0622_ clknet_leaf_97_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[1\]\[22\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_95_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5731_ _2819_ _0508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5662_ _0920_ _2778_ _2782_ _0476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_30_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4613_ soc.spi_video_ram_1.write_fifo.fifo_mem\[4\]\[2\] soc.spi_video_ram_1.fifo_in_data\[2\]
+ _2058_ _2061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5593_ soc.spi_video_ram_1.fifo_in_address\[12\] soc.spi_video_ram_1.write_fifo.fifo_mem\[5\]\[28\]
+ _2704_ _2737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_30_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4544_ _2022_ _2023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_144_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6214_ _0089_ clknet_leaf_143_wb_clk_i soc.spi_video_ram_1.state_counter\[9\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4475_ soc.video_generator_1.v_count\[0\] _1458_ _1980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_3426_ _0907_ soc.cpu.AReg.data\[9\] _1012_ soc.ram_data_out\[9\] _1030_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6145_ _0025_ clknet_leaf_67_wb_clk_i soc.ram_encoder_0.output_buffer\[6\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3357_ _0963_ _0964_ _0965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_85_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6076_ soc.spi_video_ram_1.write_fifo.fifo_mem\[2\]\[11\] soc.spi_video_ram_1.fifo_in_data\[11\]
+ _3031_ _3033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5027_ _2330_ _2332_ _2336_ _2340_ _2341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3288_ _0886_ _0899_ _0875_ _0900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_39_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_73_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_26_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1906 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_130_wb_clk_i clknet_4_2_0_wb_clk_i clknet_leaf_130_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_1939 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1928 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1917 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6978_ net57 net56 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_142_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5929_ _2954_ _0571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_139_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_72_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4260_ _1584_ _1790_ _1791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_79_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3211_ _0757_ _0802_ _0824_ _0825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4191_ _1581_ _1726_ _1727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_95_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3142_ _0749_ _0751_ _0755_ _0756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_10_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3073_ soc.spi_video_ram_1.write_fifo.write_pointer\[0\] _0693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_82_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3975_ soc.ram_encoder_0.output_buffer\[11\] _1527_ _1542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_51_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6763_ _0605_ clknet_leaf_126_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[1\]\[5\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6694_ _0536_ clknet_leaf_50_wb_clk_i soc.synch_hack_writeM vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5714_ soc.spi_video_ram_1.write_fifo.fifo_mem\[6\]\[10\] soc.spi_video_ram_1.fifo_in_data\[10\]
+ _2810_ _2811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_50_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5645_ _2745_ _2770_ _2771_ _0469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_108_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5576_ _1940_ _2708_ _2728_ _0444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_117_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4527_ _0009_ _1024_ _2013_ _0109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4458_ soc.spi_video_ram_1.state_counter\[5\] _1967_ _1969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_131_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3409_ _1011_ _1013_ _1014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_77_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6128_ _1123_ _2896_ _3051_ _2572_ _0672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_98_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4389_ _1912_ _0072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6059_ soc.spi_video_ram_1.write_fifo.fifo_mem\[2\]\[3\] soc.spi_video_ram_1.fifo_in_data\[3\]
+ _3020_ _3024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_2415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1714 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1725 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1747 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1736 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1769 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_6_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3760_ _1138_ _1344_ _1348_ _1357_ _1358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_32_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5430_ _2507_ _2624_ _2625_ _2629_ _2630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_3691_ _1241_ _1288_ _1289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_126_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5361_ soc.ram_encoder_0.address\[3\] soc.ram_encoder_0.request_address\[3\] _2566_
+ _2579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_58_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5292_ _1493_ soc.ram_encoder_0.current_state\[1\] _1488_ _2530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_99_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4312_ _1839_ _0068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_114_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4243_ soc.spi_video_ram_1.write_fifo.fifo_mem\[1\]\[7\] _1775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_101_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4174_ _1595_ soc.spi_video_ram_1.write_fifo.fifo_mem\[6\]\[1\] _1709_ _1711_ _1712_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_56_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3125_ _0695_ _0699_ _0739_ _0696_ _0740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_83_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3056_ soc.spi_video_ram_1.state_counter\[9\] soc.spi_video_ram_1.state_counter\[8\]
+ soc.spi_video_ram_1.state_counter\[10\] _0677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_82_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_36_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6815_ _0657_ clknet_leaf_110_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[2\]\[28\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_23_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6746_ _0588_ clknet_leaf_74_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[0\]\[17\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_51_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3958_ _1510_ _1526_ _1528_ _0026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_109_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6677_ _0519_ clknet_leaf_37_wb_clk_i soc.cpu.AReg.clk vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3889_ _1190_ _1466_ _1462_ _1468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_136_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5628_ soc.rom_loader.current_address\[7\] _2759_ _2745_ _2760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5559_ soc.spi_video_ram_1.fifo_in_data\[11\] soc.spi_video_ram_1.write_fifo.fifo_mem\[5\]\[11\]
+ _2719_ _2720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_101_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_26_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_14_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4930_ _2274_ _0252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_64_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4861_ _1426_ _2221_ _2222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_33_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6600_ _0457_ clknet_leaf_29_wb_clk_i soc.rom_loader.current_address\[0\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_61_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3812_ _0720_ _0843_ _1402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_4792_ _2180_ _0704_ _0721_ _0703_ _1575_ _2181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_6531_ _0404_ clknet_leaf_57_wb_clk_i soc.ram_data_out\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_20_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3743_ _1326_ _1330_ _1332_ _1340_ _1341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_118_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6462_ _0335_ clknet_leaf_6_wb_clk_i soc.rom_encoder_0.current_state\[0\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3674_ _1241_ _1221_ _1272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_5413_ soc.ram_encoder_0.request_data_out\[2\] _2606_ _2616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6393_ _0266_ clknet_leaf_11_wb_clk_i soc.rom_encoder_0.request_data_out\[14\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_115_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5344_ soc.ram_encoder_0.request_data_out\[12\] _2566_ _2569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_142_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5275_ soc.ram_encoder_0.input_buffer\[2\] _2505_ _2508_ _2519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_141_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4226_ _1756_ soc.spi_video_ram_1.write_fifo.fifo_mem\[6\]\[6\] _1758_ _1759_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4157_ _1693_ _1695_ _1696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_55_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3108_ soc.spi_video_ram_1.initialized _0727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4088_ _1637_ _1640_ _1641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_leaf_37_wb_clk_i clknet_4_7_0_wb_clk_i clknet_leaf_37_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_83_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6729_ _0571_ clknet_leaf_10_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[0\]\[0\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_137_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2042 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2031 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2020 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2086 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2075 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2064 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2053 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2097 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput25 la_data_in[16] net25 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_128_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xinput36 la_data_in[26] net36 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput14 io_in[30] net14 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_10_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3390_ _0887_ soc.cpu.AReg.data\[7\] _0894_ _0996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_97_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5060_ soc.spi_video_ram_1.write_fifo.fifo_mem\[3\]\[10\] soc.spi_video_ram_1.fifo_in_data\[10\]
+ _2357_ _2360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4011_ _1522_ _1569_ _1570_ _0037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_84_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5962_ _2971_ _0587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_19_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4913_ soc.rom_encoder_0.input_buffer\[9\] _2262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_52_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5893_ net19 _2930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4844_ soc.spi_video_ram_1.fifo_write_request _2211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_60_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4775_ soc.rom_encoder_0.output_buffer\[17\] _2138_ _2167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6514_ _0387_ clknet_leaf_66_wb_clk_i soc.ram_encoder_0.request_address\[11\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3726_ _1238_ _1322_ _1323_ _1324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_119_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6445_ _0318_ clknet_leaf_51_wb_clk_i soc.cpu.DMuxJMP.sel\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3657_ _1247_ _1248_ _1251_ _1255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_6376_ _0249_ clknet_leaf_17_wb_clk_i soc.rom_encoder_0.input_buffer\[10\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3588_ _1184_ _1185_ _1182_ _1186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_114_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5327_ soc.ram_encoder_0.data_out\[7\] _2557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_88_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5258_ soc.ram_encoder_0.input_buffer\[1\] _2507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_102_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4209_ soc.spi_video_ram_1.write_fifo.fifo_mem\[7\]\[5\] _1743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5189_ _1410_ _2385_ _2452_ _2453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_84_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_16_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_25_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_26_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1171 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4560_ _1757_ _2025_ _2032_ _0123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_144_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3511_ _0904_ soc.cpu.ALU.x\[14\] _1110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4491_ _1167_ _1991_ _1992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3442_ _0926_ _1044_ _1045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_6230_ _0105_ clknet_leaf_15_wb_clk_i soc.spi_video_ram_1.fifo_in_data\[4\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_3373_ _0952_ _0980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6161_ _0041_ clknet_leaf_117_wb_clk_i soc.spi_video_ram_1.output_buffer\[2\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_40_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5112_ _2391_ _2392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_85_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6092_ soc.spi_video_ram_1.write_fifo.fifo_mem\[2\]\[19\] soc.spi_video_ram_1.fifo_in_address\[3\]
+ _3031_ _3041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_111_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5043_ soc.spi_video_ram_1.write_fifo.fifo_mem\[3\]\[2\] soc.spi_video_ram_1.fifo_in_data\[2\]
+ _2217_ _2351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5945_ _2962_ _0579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5876_ _2898_ soc.hack_clk_strobe _2919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_80_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4827_ soc.spi_video_ram_1.fifo_in_address\[8\] soc.cpu.AReg.data\[8\] _0748_ _2201_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_33_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4758_ soc.rom_encoder_0.request_address\[13\] _1650_ _2125_ soc.rom_encoder_0.output_buffer\[10\]
+ _2152_ _2153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_4689_ soc.spi_video_ram_1.state_sram_clk_counter\[4\] _2102_ _2096_ _2105_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_4_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3709_ _1216_ soc.video_generator_1.h_count\[2\] _1218_ _1307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_49_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6428_ _0301_ clknet_leaf_99_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[3\]\[14\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_134_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6359_ _0232_ clknet_leaf_127_wb_clk_i soc.spi_video_ram_1.write_fifo.write_pointer\[2\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_4
XFILLER_76_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_52_wb_clk_i clknet_4_6_0_wb_clk_i clknet_leaf_52_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_57_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_44_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_33_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3991_ soc.ram_encoder_0.output_buffer\[15\] _1527_ _1554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_62_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5730_ soc.spi_video_ram_1.write_fifo.fifo_mem\[6\]\[18\] soc.spi_video_ram_1.fifo_in_address\[2\]
+ _2810_ _2819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_15_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5661_ soc.cpu.ALU.x\[2\] _2779_ _2782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_30_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4612_ _2060_ _0147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5592_ _2736_ _0452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_128_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4543_ soc.spi_video_ram_1.write_fifo.write_pointer\[2\] _0694_ _0698_ _2022_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_144_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4474_ _1961_ _1979_ _0090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6213_ _0088_ clknet_leaf_140_wb_clk_i soc.spi_video_ram_1.state_counter\[8\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3425_ _0849_ _1028_ _1029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_6144_ _0024_ clknet_leaf_66_wb_clk_i soc.ram_encoder_0.output_buffer\[5\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3356_ _0887_ soc.cpu.AReg.data\[5\] _0894_ _0964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_58_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3287_ _0853_ _0895_ _0899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_6075_ _3032_ _0639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5026_ soc.ram_encoder_0.output_buffer\[16\] _2337_ _2338_ _2339_ _2340_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_57_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1907 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1929 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1918 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6977_ net57 net55 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_14_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5928_ soc.spi_video_ram_1.write_fifo.fifo_mem\[0\]\[0\] soc.spi_video_ram_1.fifo_in_data\[0\]
+ _2953_ _2954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_80_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5859_ _2911_ _0544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_21_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_77_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_130_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_45_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4190_ _1725_ _1726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3210_ _0783_ soc.spi_video_ram_1.output_buffer\[17\] _0824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_122_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3141_ _0751_ _0754_ _0755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_95_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3072_ _0687_ _0692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_36_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6831_ _0673_ clknet_leaf_48_wb_clk_i soc.ram_encoder_0.data_out\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_51_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3974_ soc.ram_encoder_0.output_buffer\[7\] _1520_ _1530_ soc.ram_encoder_0.request_data_out\[3\]
+ _1540_ _1541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_6762_ _0604_ clknet_leaf_130_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[1\]\[4\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6693_ _0535_ clknet_leaf_37_wb_clk_i soc.hack_clk_strobe vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5713_ _2797_ _2810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_5644_ soc.rom_loader.current_address\[12\] _2769_ _2771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_31_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5575_ soc.spi_video_ram_1.fifo_in_address\[3\] _2705_ _2728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xclkbuf_4_3_0_wb_clk_i clknet_0_wb_clk_i clknet_4_3_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_132_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4526_ soc.spi_video_ram_1.fifo_in_data\[8\] _2007_ _2013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4457_ _1961_ _1967_ _1968_ _0084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_3408_ _0907_ soc.cpu.AReg.data\[8\] _1012_ soc.ram_data_out\[8\] _1013_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6127_ _1108_ _2896_ _3051_ _2570_ _0671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_59_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4388_ soc.spi_video_ram_1.output_buffer\[8\] _1612_ _1825_ _1911_ _1912_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_112_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3339_ soc.ram_data_out\[4\] _0869_ _0868_ net41 _0854_ _0948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_86_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6058_ _3023_ _0631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_22_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5009_ _2325_ _0280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_26_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1715 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1704 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1748 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1737 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1726 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1759 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_20_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3690_ _1278_ _1287_ _1288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_127_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_126_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5360_ _2578_ _0378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_141_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5291_ _2528_ _2505_ _2529_ _0358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4311_ soc.spi_video_ram_1.output_buffer\[12\] _1612_ _1825_ _1838_ _1839_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_114_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_102_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4242_ soc.spi_video_ram_1.write_fifo.fifo_mem\[2\]\[7\] soc.spi_video_ram_1.write_fifo.fifo_mem\[3\]\[7\]
+ _1600_ _1774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_68_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4173_ _1710_ _1711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_83_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_109_wb_clk_i clknet_4_10_0_wb_clk_i clknet_leaf_109_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_3124_ _0701_ _0738_ _0739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_49_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3055_ _0675_ _0676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_82_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_70_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6814_ _0656_ clknet_leaf_99_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[2\]\[27\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3957_ soc.ram_encoder_0.output_buffer\[7\] _1527_ _1528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6745_ _0587_ clknet_leaf_79_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[0\]\[16\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_23_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6676_ _0518_ clknet_leaf_116_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[6\]\[28\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3888_ _1460_ _1466_ _1467_ _0017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_118_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5627_ _2746_ _2758_ _2759_ _0463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_117_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5558_ _2704_ _2719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_133_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4509_ soc.spi_video_ram_1.fifo_in_data\[0\] _2003_ _2004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_120_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5489_ _0676_ _2674_ _0411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_78_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_27_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_2279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_127_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_68_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_7_wb_clk_i clknet_4_1_0_wb_clk_i clknet_leaf_7_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_2_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4860_ soc.rom_encoder_0.current_state\[1\] _1406_ _2221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_60_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3811_ _1388_ _1399_ _1401_ _0720_ net72 vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
X_6530_ _0403_ clknet_leaf_57_wb_clk_i soc.ram_data_out\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4791_ soc.spi_video_ram_1.state_sram_clk_counter\[0\] _0684_ _0715_ _2180_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_20_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_32_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_9_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3742_ _1243_ _1335_ _1339_ _1340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_6461_ _0334_ clknet_leaf_7_wb_clk_i soc.rom_encoder_0.sram_sio_oe vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3673_ _1261_ _1270_ _1265_ _1271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5412_ _0689_ _2615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_6392_ _0265_ clknet_leaf_37_wb_clk_i soc.rom_encoder_0.request_data_out\[13\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5343_ soc.ram_encoder_0.data_out\[12\] _2568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5274_ soc.ram_encoder_0.input_buffer\[6\] _2518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_102_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4225_ _1724_ _1757_ _1758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_68_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4156_ soc.spi_video_ram_1.current_state\[4\] _1694_ _1695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_83_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_56_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3107_ soc.spi_video_ram_1.current_state\[3\] _0725_ _0726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_28_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4087_ soc.ram_encoder_0.output_bits_left\[2\] soc.ram_encoder_0.output_bits_left\[3\]
+ _1640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_56_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_70_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_77_wb_clk_i clknet_4_12_0_wb_clk_i clknet_leaf_77_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_4989_ _2293_ _2310_ _2311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_51_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6728_ _0570_ net87 soc.gpio_i_stored\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_109_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6659_ _0501_ clknet_leaf_92_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[6\]\[11\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_20_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2010 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2043 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2032 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2021 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2076 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2065 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2054 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2098 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2087 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput15 io_in[31] net15 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput37 la_data_in[28] net37 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput26 la_data_in[17] net26 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_7_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_97_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4010_ soc.ram_encoder_0.output_buffer\[18\] _1509_ _1570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_96_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_38_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5961_ soc.spi_video_ram_1.write_fifo.fifo_mem\[0\]\[16\] soc.spi_video_ram_1.fifo_in_address\[0\]
+ _2964_ _2971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_65_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4912_ _2260_ _2242_ _2261_ _0247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_34_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5892_ net85 soc.hack_clk_strobe _2929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_34_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4843_ _0727_ _0722_ _0691_ _0229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_33_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4774_ soc.rom_encoder_0.output_buffer\[13\] _2163_ _2165_ _1435_ _1441_ _2166_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_6513_ _0386_ clknet_4_13_0_wb_clk_i soc.ram_encoder_0.request_address\[10\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3725_ _1311_ _1264_ _1323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_20_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6444_ _0317_ clknet_leaf_16_wb_clk_i soc.cpu.DMuxJMP.sel\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_134_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3656_ _1202_ _1206_ _1234_ _1201_ _1253_ _1254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
X_6375_ _0248_ clknet_leaf_21_wb_clk_i soc.rom_encoder_0.input_buffer\[9\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3587_ _1180_ _1183_ _1171_ _1185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5326_ _2555_ _2542_ _2556_ _0366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_103_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xclkbuf_leaf_124_wb_clk_i clknet_4_3_0_wb_clk_i clknet_leaf_124_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_130_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5257_ _2502_ _2504_ _2506_ _0347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_88_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4208_ _1595_ soc.spi_video_ram_1.write_fifo.fifo_mem\[4\]\[5\] _1741_ _1742_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5188_ _1426_ _1408_ _1419_ _1425_ _2452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4139_ _1522_ _1679_ _1680_ _0054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_110_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_106_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_35_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3510_ _0883_ _1108_ _1109_ soc.cpu.PC.in\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4490_ _1984_ _1990_ _1991_ _0094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_144_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3441_ _1011_ _1043_ _1044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_6_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3372_ _0974_ _0978_ _0979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_6160_ _0040_ clknet_leaf_117_wb_clk_i soc.spi_video_ram_1.output_buffer\[3\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5111_ _1407_ soc.rom_encoder_0.current_state\[1\] _2390_ _2391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_33_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6091_ _3040_ _0647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5042_ _2350_ _0288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_81_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_19_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5944_ soc.spi_video_ram_1.write_fifo.fifo_mem\[0\]\[8\] soc.spi_video_ram_1.fifo_in_data\[8\]
+ _2953_ _2962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_41_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5875_ _2897_ _0553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4826_ _2200_ _0222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_22_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4757_ soc.rom_encoder_0.request_data_out\[6\] _1481_ _2152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_21_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4688_ soc.spi_video_ram_1.state_sram_clk_counter\[4\] _2102_ _2104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_3708_ _1260_ _1301_ _1287_ _1265_ _1306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_108_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3639_ _1230_ _1232_ _1233_ _1237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_6427_ _0300_ clknet_leaf_108_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[3\]\[13\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_122_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6358_ _0231_ clknet_leaf_130_wb_clk_i soc.spi_video_ram_1.write_fifo.write_pointer\[1\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5309_ _2537_ _2545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_88_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6289_ _0164_ clknet_leaf_82_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[4\]\[18\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_112_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_92_wb_clk_i clknet_4_11_0_wb_clk_i clknet_leaf_92_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_17_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xclkbuf_leaf_21_wb_clk_i clknet_4_4_0_wb_clk_i clknet_leaf_21_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_72_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_32_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3990_ soc.ram_encoder_0.request_address\[14\] _1514_ _1530_ soc.ram_encoder_0.request_data_out\[7\]
+ _1552_ _1553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_23_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5660_ _0902_ _2778_ _2781_ _0475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_15_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4611_ soc.spi_video_ram_1.write_fifo.fifo_mem\[4\]\[1\] soc.spi_video_ram_1.fifo_in_data\[1\]
+ _2058_ _2060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_129_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5591_ soc.spi_video_ram_1.fifo_in_address\[11\] soc.spi_video_ram_1.write_fifo.fifo_mem\[5\]\[27\]
+ _2719_ _2736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4542_ _2003_ _1669_ _2021_ _0116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_8_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4473_ soc.spi_video_ram_1.state_counter\[10\] _1978_ _1979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_116_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3424_ _0850_ soc.cpu.ALU.x\[9\] _1028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6212_ _0087_ clknet_leaf_143_wb_clk_i soc.spi_video_ram_1.state_counter\[7\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_144_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3355_ soc.ram_data_out\[5\] _0869_ _0868_ net42 _0907_ _0963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XTAP_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6143_ _0023_ clknet_leaf_1_wb_clk_i net64 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3286_ soc.cpu.ALU.f _0897_ _0898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6074_ soc.spi_video_ram_1.write_fifo.fifo_mem\[2\]\[10\] soc.spi_video_ram_1.fifo_in_data\[10\]
+ _3031_ _3032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_58_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5025_ _1492_ _1494_ _2339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_100_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1908 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6976_ net57 net54 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_13_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5927_ _2952_ _2953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_5858_ soc.ram_encoder_0.address\[7\] soc.cpu.AReg.data\[7\] _2902_ _2911_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_16_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5789_ _2531_ _2861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_4809_ _1796_ _2192_ _0213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_119_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_71_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_69_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_140_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3140_ soc.spi_video_ram_1.buffer_index\[4\] _0753_ _0754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_67_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3071_ _0690_ _0691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_54_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6830_ _0672_ clknet_leaf_50_wb_clk_i soc.ram_encoder_0.data_out\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_36_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6761_ _0603_ clknet_leaf_10_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[1\]\[3\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3973_ soc.ram_encoder_0.request_address\[10\] _1513_ _1540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_5712_ _2809_ _0499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_50_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6692_ _0534_ net86 soc.cpu.PC.REG.data\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5643_ soc.rom_loader.current_address\[12\] _2769_ _2770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_117_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5574_ _1615_ _2707_ _2727_ _0443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_102_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4525_ _0009_ _1002_ _2012_ _0108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_144_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_117_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4456_ soc.spi_video_ram_1.state_counter\[4\] _1965_ _1968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_132_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3407_ _0854_ _0858_ _1012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_4387_ _1821_ _1904_ _1909_ _1850_ _1910_ _1911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_6126_ _1092_ _2896_ _3051_ _2568_ _0670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_3338_ _0849_ _0946_ _0947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3269_ _0846_ _0847_ _0848_ _0878_ _0881_ _0855_ soc.cpu.PC.in\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__oai222_2
XFILLER_22_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6057_ soc.spi_video_ram_1.write_fifo.fifo_mem\[2\]\[2\] soc.spi_video_ram_1.fifo_in_data\[2\]
+ _3020_ _3023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_2417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5008_ _2324_ soc.rom_encoder_0.request_address\[12\] _2271_ _2325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_39_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1705 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1749 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1716 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1727 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_89_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_45_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5290_ soc.ram_encoder_0.input_buffer\[7\] _2503_ _0675_ _2529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4310_ _1821_ _1830_ _1834_ _1837_ _1838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_4241_ _1592_ _1769_ _1772_ _1605_ _1773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_141_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4172_ _1586_ _1710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_67_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3123_ _0694_ soc.spi_video_ram_1.write_fifo.write_pointer\[0\] _0738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_55_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3054_ _0674_ _0675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_82_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6813_ _0655_ clknet_leaf_99_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[2\]\[26\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3956_ _1509_ _1527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_6744_ _0586_ clknet_leaf_73_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[0\]\[15\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_23_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6675_ _0517_ clknet_leaf_97_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[6\]\[27\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5626_ soc.rom_loader.current_address\[6\] _2757_ _2759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_31_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3887_ soc.video_generator_1.h_count\[4\] _1464_ _1467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5557_ _2718_ _0435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_144_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5488_ soc.ram_encoder_0.current_state\[1\] _2670_ _2671_ _1557_ _2674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_4508_ _0748_ _2003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_144_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4439_ soc.spi_video_ram_1.write_fifo.read_pointer\[2\] _1954_ _1956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_133_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6109_ _3049_ _0656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_74_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_30_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_23_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_10_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_49_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3810_ _0764_ _0770_ _1400_ _1401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4790_ _0776_ _2177_ _2179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_33_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3741_ _1140_ _1338_ _1199_ _1339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_119_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6460_ _0333_ clknet_leaf_7_wb_clk_i net62 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3672_ _1217_ _1269_ _1270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_5411_ _2436_ _2614_ _0393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6391_ _0264_ clknet_leaf_32_wb_clk_i soc.rom_encoder_0.request_data_out\[12\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_63_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5342_ _2565_ _2538_ _2567_ _0371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_114_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5273_ _2516_ _2504_ _2517_ _0352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_115_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4224_ soc.spi_video_ram_1.write_fifo.fifo_mem\[7\]\[6\] _1757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_68_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4155_ _0681_ _1607_ _1694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_110_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3106_ soc.spi_video_ram_1.state_sram_clk_counter\[2\] _0713_ _0725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_4086_ _1635_ _1638_ _1639_ _0042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_83_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4988_ soc.cpu.PC.REG.data\[7\] _2310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3939_ soc.ram_encoder_0.current_state\[1\] _1502_ _1512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6727_ _0569_ net91 soc.gpio_i_stored\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_127_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6658_ _0500_ clknet_leaf_90_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[6\]\[10\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_125_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_46_wb_clk_i clknet_4_6_0_wb_clk_i clknet_leaf_46_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_5609_ _2744_ _2746_ _2747_ _0457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_105_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6589_ net26 clknet_leaf_94_wb_clk_i soc.rom_encoder_0.data_out\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_105_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2000 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2033 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2022 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2011 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2077 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2066 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2055 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2044 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2099 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2088 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_11_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput27 la_data_in[18] net27 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_11_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput16 io_in[32] net16 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput38 la_data_in[2] net38 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_6_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_115_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_2_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5960_ _2970_ _0586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4911_ soc.rom_encoder_0.input_buffer\[4\] _2241_ _2250_ _2261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5891_ _2471_ _2928_ _0559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_45_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4842_ _0691_ _2210_ _0228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4773_ soc.rom_encoder_0.current_state\[1\] _2164_ _2165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6512_ _0385_ clknet_leaf_64_wb_clk_i soc.ram_encoder_0.request_address\[9\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3724_ _1309_ _1321_ _1239_ _1322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_107_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6443_ _0316_ clknet_leaf_7_wb_clk_i soc.rom_encoder_0.initialized vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3655_ _1176_ _1186_ _1253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_6374_ _0247_ clknet_leaf_18_wb_clk_i soc.rom_encoder_0.input_buffer\[8\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3586_ _1180_ _1183_ _1184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_5325_ soc.ram_encoder_0.request_data_out\[6\] _2545_ _2556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5256_ net1 _2505_ _2250_ _2506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_88_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4207_ _1596_ _1740_ _1741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5187_ _2436_ _2451_ _0332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4138_ soc.ram_encoder_0.output_buffer\[3\] _1509_ _1680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_83_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4069_ soc.spi_video_ram_1.write_fifo.fifo_mem\[0\]\[17\] soc.spi_video_ram_1.write_fifo.fifo_mem\[1\]\[17\]
+ soc.spi_video_ram_1.write_fifo.fifo_mem\[2\]\[17\] soc.spi_video_ram_1.write_fifo.fifo_mem\[3\]\[17\]
+ _1585_ _1588_ _1624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_58_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_25_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_79_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_8_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3440_ _0907_ soc.cpu.AReg.data\[10\] _1012_ soc.ram_data_out\[10\] _1043_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3371_ _0853_ _0977_ _0978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_112_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6090_ soc.spi_video_ram_1.write_fifo.fifo_mem\[2\]\[18\] soc.spi_video_ram_1.fifo_in_address\[2\]
+ _3031_ _3040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5110_ _1403_ _2389_ _2390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5041_ soc.spi_video_ram_1.write_fifo.fifo_mem\[3\]\[1\] soc.spi_video_ram_1.fifo_in_data\[1\]
+ _2217_ _2350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_38_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_0_wb_clk_i wb_clk_i clknet_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_92_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5943_ _2961_ _0578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5874_ _2899_ _0552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_80_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4825_ soc.spi_video_ram_1.fifo_in_address\[7\] soc.cpu.AReg.data\[7\] _0748_ _2200_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_61_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4756_ _2122_ _2150_ _2151_ _0201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_134_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4687_ _2102_ _2103_ _0179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3707_ _1271_ _1304_ _1305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6426_ _0299_ clknet_leaf_74_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[3\]\[12\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3638_ _1202_ _1235_ _1236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_3569_ soc.video_generator_1.v_count\[4\] _1167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
X_6357_ _0230_ clknet_leaf_130_wb_clk_i soc.spi_video_ram_1.write_fifo.write_pointer\[0\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_103_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5308_ soc.ram_encoder_0.data_out\[1\] _2544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_103_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6288_ _0163_ clknet_leaf_85_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[4\]\[17\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5239_ soc.ram_encoder_0.toggled_sram_sck _2491_ _2492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_48_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_84_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_72_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xclkbuf_leaf_61_wb_clk_i clknet_4_13_0_wb_clk_i clknet_leaf_61_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XPHY_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_130_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_12_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_137_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_47_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4610_ _2059_ _0146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_30_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5590_ _2735_ _0451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4541_ soc.spi_video_ram_1.fifo_in_data\[15\] _2018_ _2021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_144_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4472_ soc.spi_video_ram_1.state_counter\[9\] _1975_ _1978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_144_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3423_ _1005_ _1008_ _1016_ _1027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6211_ _0086_ clknet_leaf_143_wb_clk_i soc.spi_video_ram_1.state_counter\[6\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6142_ _0022_ clknet_leaf_0_wb_clk_i soc.video_generator_1.h_count\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_135_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3354_ _0923_ _0961_ _0962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3285_ _0877_ _0896_ _0897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_6073_ _3018_ _3031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XTAP_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5024_ soc.ram_encoder_0.initializing_step\[1\] soc.ram_encoder_0.initializing_step\[0\]
+ _2331_ soc.ram_encoder_0.initializing_step\[2\] _2338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6975_ net53 net52 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1909 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5926_ _2951_ _2952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_139_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5857_ _2910_ _0543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_10_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5788_ soc.cpu.PC.REG.data\[4\] _2859_ _2860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_4808_ soc.spi_video_ram_1.buffer_index\[5\] _2191_ _2192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_21_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4739_ soc.rom_encoder_0.output_buffer\[9\] _2138_ _2139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_135_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6409_ _0282_ clknet_leaf_23_wb_clk_i soc.rom_encoder_0.request_address\[14\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_131_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_40_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3070_ _0689_ _0690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_79_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_63_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6760_ _0602_ clknet_leaf_10_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[1\]\[2\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_23_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3972_ _1510_ _1538_ _1539_ _0029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_93_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5711_ soc.spi_video_ram_1.write_fifo.fifo_mem\[6\]\[9\] soc.spi_video_ram_1.fifo_in_data\[9\]
+ _2799_ _2809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_51_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6691_ _0533_ net86 soc.cpu.PC.REG.data\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5642_ _2745_ _2768_ _2769_ _0468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_31_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5573_ soc.spi_video_ram_1.fifo_in_address\[2\] _2705_ _2727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_144_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4524_ soc.spi_video_ram_1.fifo_in_data\[7\] _2007_ _2012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_144_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4455_ soc.spi_video_ram_1.state_counter\[4\] _1965_ _1967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_3406_ soc.cpu.ALU.zy _1011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_4386_ soc.video_generator_1.v_count\[2\] _1129_ _0729_ _1910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6125_ _1069_ _2896_ _3051_ _2565_ _0669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_98_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3337_ _0850_ soc.cpu.ALU.x\[4\] _0946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3268_ _0880_ _0881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6056_ _3022_ _0630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5007_ soc.cpu.PC.REG.data\[12\] soc.rom_loader.current_address\[12\] _2292_ _2324_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3199_ _0808_ _0809_ _0811_ _0812_ _0813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_26_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1739 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1717 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1728 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5909_ net80 _2936_ _2861_ _2940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_22_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_22_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_60_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_5_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4240_ _1595_ soc.spi_video_ram_1.write_fifo.fifo_mem\[6\]\[7\] _1771_ _1711_ _1772_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_4171_ _1585_ _1708_ _1709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_45_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3122_ _0735_ _0737_ _0691_ _0004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_82_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3053_ net18 _0674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_4
XFILLER_64_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6812_ _0654_ clknet_leaf_111_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[2\]\[25\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_36_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3955_ soc.ram_encoder_0.request_address\[6\] _1514_ _1520_ soc.ram_encoder_0.output_buffer\[3\]
+ _1526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6743_ _0585_ clknet_leaf_98_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[0\]\[14\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6674_ _0516_ clknet_leaf_101_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[6\]\[26\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_32_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5625_ soc.rom_loader.current_address\[6\] _2757_ _2758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3886_ soc.video_generator_1.h_count\[4\] _1464_ _1466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
Xclkbuf_leaf_118_wb_clk_i clknet_4_9_0_wb_clk_i clknet_leaf_118_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_5556_ soc.spi_video_ram_1.fifo_in_data\[10\] soc.spi_video_ram_1.write_fifo.fifo_mem\[5\]\[10\]
+ _2705_ _2718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_3_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5487_ _2672_ _2673_ _0410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4507_ _1142_ _2001_ _2002_ _1984_ _0100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_132_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4438_ _0675_ _1955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_101_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4369_ _1584_ soc.spi_video_ram_1.write_fifo.fifo_mem\[6\]\[14\] _1893_ _1590_ _1894_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_101_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6108_ soc.spi_video_ram_1.write_fifo.fifo_mem\[2\]\[27\] soc.spi_video_ram_1.fifo_in_address\[11\]
+ _3019_ _3049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_132_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6039_ _3012_ _0623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_10_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_20_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3740_ soc.video_generator_1.v_count\[1\] _1168_ _1129_ _1337_ _1338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_12_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3671_ _1268_ _1219_ _1220_ _1269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6390_ _0263_ clknet_leaf_37_wb_clk_i soc.rom_encoder_0.request_data_out\[11\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5410_ soc.ram_data_out\[1\] _2603_ _2613_ _2614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_12_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5341_ soc.ram_encoder_0.request_data_out\[11\] _2566_ _2567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_56_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5272_ soc.ram_encoder_0.input_buffer\[1\] _2505_ _2508_ _2517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_141_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4223_ _1755_ _1756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_95_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4154_ _1352_ _1353_ _1354_ _1693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_4085_ _1497_ _1635_ soc.ram_encoder_0.output_bits_left\[4\] _1639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_110_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_83_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3105_ _0691_ _0724_ _0005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_83_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6726_ _0568_ net87 soc.gpio_i_stored\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4987_ _2309_ _0274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3938_ soc.ram_encoder_0.output_bits_left\[4\] _1498_ _1511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_6657_ _0499_ clknet_leaf_80_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[6\]\[9\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_20_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3869_ net67 _1432_ _1454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6588_ net25 clknet_leaf_33_wb_clk_i soc.rom_encoder_0.data_out\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5608_ soc.rom_loader.current_address\[0\] _0473_ _2747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5539_ _1705_ _2707_ _2709_ _0426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_117_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_86_wb_clk_i clknet_4_9_0_wb_clk_i clknet_leaf_86_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_2_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_leaf_15_wb_clk_i clknet_4_6_0_wb_clk_i clknet_leaf_15_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_47_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2001 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2034 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2023 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2012 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2067 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2056 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2045 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2089 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2078 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput17 io_in[33] net17 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_122_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput28 la_data_in[19] net28 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput39 la_data_in[3] net39 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_108_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_92_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4910_ soc.rom_encoder_0.input_buffer\[8\] _2260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_19_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5890_ soc.boot_loading_offset\[4\] _2927_ _2928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4841_ soc.spi_video_ram_1.start_read _0705_ _2209_ _2210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_45_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4772_ soc.rom_encoder_0.request_data_out\[9\] _1434_ _2164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6511_ _0384_ clknet_leaf_65_wb_clk_i soc.ram_encoder_0.request_address\[8\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3723_ _1306_ _1319_ _1320_ _1321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3654_ _1247_ _1248_ _1251_ _1252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6442_ _0315_ clknet_leaf_110_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[3\]\[28\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_127_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_115_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6373_ _0246_ clknet_leaf_16_wb_clk_i soc.rom_encoder_0.input_buffer\[7\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3585_ soc.boot_loading_offset\[4\] _1182_ _1183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_138_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_103_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5324_ soc.ram_encoder_0.data_out\[6\] _2555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_88_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5255_ _2503_ _2505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_88_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4206_ soc.spi_video_ram_1.write_fifo.fifo_mem\[5\]\[5\] _1740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_111_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5186_ _0846_ _2393_ _2450_ _2451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_68_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4137_ soc.ram_encoder_0.request_address\[2\] _1514_ _1679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_84_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4068_ _1578_ _1622_ _1623_ _0040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_25_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_133_wb_clk_i clknet_4_2_0_wb_clk_i clknet_leaf_133_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_12_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6709_ _0551_ clknet_leaf_56_wb_clk_i soc.ram_encoder_0.address\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_20_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_79_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_19_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_16_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3370_ _0975_ _0976_ _0977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_111_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5040_ _2349_ _0287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_2_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5942_ soc.spi_video_ram_1.write_fifo.fifo_mem\[0\]\[7\] soc.spi_video_ram_1.fifo_in_data\[7\]
+ _2953_ _2961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5873_ _2918_ _0551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_80_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_22_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4824_ _2199_ _0221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_33_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4755_ soc.rom_encoder_0.output_buffer\[13\] _2138_ _2151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3706_ _1286_ _1261_ _1303_ _1304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4686_ soc.spi_video_ram_1.state_sram_clk_counter\[3\] _2100_ _2096_ _2103_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6425_ _0298_ clknet_leaf_92_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[3\]\[11\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3637_ _1206_ _1234_ _1235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_143_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3568_ _1163_ _1165_ _1166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_6356_ _0229_ clknet_leaf_134_wb_clk_i soc.spi_video_ram_1.initialized vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5307_ _2541_ _2542_ _2543_ _0360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_89_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3499_ _0926_ _1098_ _1099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_6287_ _0162_ clknet_leaf_121_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[4\]\[16\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5238_ soc.ram_encoder_0.request_write _1511_ _2490_ _2491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_57_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5169_ _2258_ _2413_ _2414_ _2437_ _2438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_56_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_24_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_123_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_30_wb_clk_i clknet_4_5_0_wb_clk_i clknet_leaf_30_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_106_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_144_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4540_ _2003_ _1123_ _2020_ _0115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_144_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4471_ _1961_ _1977_ _0089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3422_ _1010_ _1015_ _1026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6210_ _0085_ clknet_leaf_139_wb_clk_i soc.spi_video_ram_1.state_counter\[5\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_48_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6141_ _0021_ clknet_leaf_0_wb_clk_i soc.video_generator_1.h_count\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_124_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_112_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3353_ _0904_ soc.cpu.ALU.x\[5\] _0961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3284_ _0853_ _0886_ _0895_ _0896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_6072_ _3030_ _0638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_58_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5023_ _1489_ _1512_ _1518_ _2337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_112_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6974_ net53 net51 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_53_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_53_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_80_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5925_ soc.spi_video_ram_1.write_fifo.write_pointer\[2\] _0694_ _0698_ _2951_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_110_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5856_ soc.ram_encoder_0.address\[6\] soc.cpu.AReg.data\[6\] _2902_ _2910_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_22_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4807_ _0749_ _0753_ _2176_ _2184_ _2191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_21_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5787_ _2300_ _2856_ _2859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4738_ _1670_ _2138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_134_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4669_ _2089_ _0689_ _2090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6408_ _0281_ clknet_leaf_21_wb_clk_i soc.rom_encoder_0.request_address\[13\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_122_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6339_ _0009_ clknet_leaf_15_wb_clk_i soc.spi_video_ram_1.fifo_write_request vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_62_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_135_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_62_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_126_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_141_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_35_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3971_ soc.ram_encoder_0.output_buffer\[10\] _1527_ _1539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_90_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5710_ _2808_ _0498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6690_ _0532_ net86 soc.cpu.PC.REG.data\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_86_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5641_ soc.rom_loader.current_address\[11\] _2767_ _2769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_5572_ _1625_ _2707_ _2726_ _0442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_116_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4523_ _0009_ _0989_ _2011_ _0107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_144_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_132_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4454_ _1961_ _1965_ _1966_ _0083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_131_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3405_ _0849_ _1009_ _1010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_4385_ _1761_ _1905_ _1908_ _1909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_113_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6124_ _1058_ _2896_ _3051_ _2563_ _0668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_86_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3336_ _0937_ _0944_ _0939_ _0945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XTAP_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6055_ soc.spi_video_ram_1.write_fifo.fifo_mem\[2\]\[1\] soc.spi_video_ram_1.fifo_in_data\[1\]
+ _3020_ _3022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3267_ soc.cpu.instruction\[15\] _0879_ _0880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_86_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5006_ _2323_ _0279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3198_ soc.spi_video_ram_1.output_buffer\[10\] soc.spi_video_ram_1.output_buffer\[11\]
+ _0757_ _0812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_2419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1718 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1729 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1707 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5908_ _0920_ _2936_ _2939_ _0565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_14_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5839_ soc.synch_hack_writeM _2899_ _2900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_108_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_6_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_92_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_45_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4170_ soc.spi_video_ram_1.write_fifo.fifo_mem\[7\]\[1\] _1708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_45_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3121_ soc.spi_video_ram_1.initialized _0008_ _0737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_55_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6811_ _0653_ clknet_leaf_108_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[2\]\[24\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_90_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3954_ _1510_ _1524_ _1525_ _0025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6742_ _0584_ clknet_leaf_109_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[0\]\[13\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_32_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6673_ _0515_ clknet_leaf_111_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[6\]\[25\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3885_ _1460_ _1464_ _1465_ _0016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_32_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5624_ _2746_ _2756_ _2757_ _0462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_118_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5555_ _1804_ _2707_ _2717_ _0434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_133_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5486_ _1488_ _2670_ _1955_ _2673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_105_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4506_ _1142_ _2001_ _2002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4437_ _1461_ _1953_ _1954_ _0078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_99_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6107_ _3048_ _0655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4368_ _1755_ _1892_ _1893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3319_ net40 _0929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_100_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4299_ soc.spi_video_ram_1.write_fifo.fifo_mem\[4\]\[11\] soc.spi_video_ram_1.write_fifo.fifo_mem\[5\]\[11\]
+ soc.spi_video_ram_1.write_fifo.fifo_mem\[6\]\[11\] soc.spi_video_ram_1.write_fifo.fifo_mem\[7\]\[11\]
+ _1583_ _1586_ _1827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6038_ soc.spi_video_ram_1.fifo_in_address\[7\] soc.spi_video_ram_1.write_fifo.fifo_mem\[1\]\[23\]
+ _2985_ _3012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_27_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_66_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_15_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_26_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_109_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_50_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_2_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_4_2_0_wb_clk_i clknet_0_wb_clk_i clknet_4_2_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_73_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_13_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3670_ soc.video_generator_1.h_count\[1\] _1216_ _1268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_115_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5340_ _2537_ _2566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_142_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5271_ soc.ram_encoder_0.input_buffer\[5\] _2516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_49_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4222_ _1582_ _1755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_68_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4153_ _0720_ _0704_ _1692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_4084_ soc.ram_encoder_0.output_bits_left\[2\] _1636_ _1637_ _1638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_96_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3104_ soc.spi_video_ram_1.current_state\[0\] _0692_ _0709_ _0723_ _0724_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_49_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4986_ _2308_ soc.rom_encoder_0.request_address\[6\] _2287_ _2309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_12_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3937_ _1509_ _1510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_6725_ _0567_ net89 soc.gpio_i_stored\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_51_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_20_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3868_ soc.rom_encoder_0.output_buffer\[19\] _1436_ _1452_ _1441_ _1453_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_20_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6656_ _0498_ clknet_leaf_120_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[6\]\[8\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6587_ net24 clknet_leaf_33_wb_clk_i soc.rom_encoder_0.data_out\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5607_ _2745_ _2746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_3799_ _1389_ _1390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5538_ soc.spi_video_ram_1.fifo_in_data\[1\] _2708_ _2709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_132_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5469_ soc.ram_encoder_0.request_data_out\[15\] _2605_ _2659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_120_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_19_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_55_wb_clk_i clknet_4_13_0_wb_clk_i clknet_leaf_55_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_2024 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2013 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2002 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2068 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2057 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2035 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2046 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2079 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xinput18 la_data_in[0] net18 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_128_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput29 la_data_in[1] net29 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xcaravel_hack_soc_220 wbs_dat_o[27] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_10_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_96_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_93_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4840_ _1356_ _1455_ _2208_ _0705_ _2209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_34_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_20_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1890 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6510_ _0383_ clknet_leaf_65_wb_clk_i soc.ram_encoder_0.request_address\[7\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4771_ _1421_ _1442_ _2163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_33_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3722_ _1261_ _1266_ _1279_ _1286_ _1320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_3653_ _1249_ _1250_ _1251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_6441_ _0314_ clknet_leaf_99_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[3\]\[27\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6372_ _0245_ clknet_leaf_17_wb_clk_i soc.rom_encoder_0.input_buffer\[6\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5323_ _2553_ _2542_ _2554_ _0365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3584_ soc.video_generator_1.v_count\[4\] _1181_ _1163_ _1182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_138_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5254_ _2503_ _2504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_102_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5185_ _2266_ _2395_ _2391_ _2449_ _2450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_4205_ _1736_ _1738_ _1739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4136_ _1522_ _1677_ _1678_ _0053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_110_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4067_ soc.spi_video_ram_1.output_buffer\[3\] _1612_ _1623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_44_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4969_ _2296_ soc.rom_encoder_0.request_address\[1\] _2287_ _2297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6708_ _0550_ clknet_leaf_53_wb_clk_i soc.ram_encoder_0.address\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_20_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6639_ _0481_ net90 soc.cpu.ALU.x\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_137_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_90_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_97_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5941_ _2960_ _0577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_19_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5872_ soc.ram_encoder_0.address\[14\] soc.cpu.AReg.data\[14\] _2902_ _2918_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_61_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_0_wb_clk_i clknet_4_0_0_wb_clk_i clknet_leaf_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_4823_ soc.spi_video_ram_1.fifo_in_address\[6\] soc.cpu.AReg.data\[6\] _2018_ _2199_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_21_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4754_ soc.rom_encoder_0.request_address\[12\] _1650_ _2125_ soc.rom_encoder_0.output_buffer\[9\]
+ _2149_ _2150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_3705_ _1280_ _1300_ _1290_ _1217_ _1302_ _1303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_119_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4685_ soc.spi_video_ram_1.state_sram_clk_counter\[3\] _2100_ _2102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_6424_ _0297_ clknet_leaf_85_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[3\]\[10\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3636_ _1203_ _1205_ _1230_ _1232_ _1233_ _1234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_108_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6355_ _0228_ clknet_leaf_132_wb_clk_i soc.spi_video_ram_1.start_read vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3567_ soc.video_generator_1.v_count\[3\] _1164_ _1143_ _1142_ _1165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
X_5306_ soc.ram_encoder_0.request_data_out\[0\] _2538_ _2543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_103_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6286_ _0161_ clknet_leaf_93_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[4\]\[15\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5237_ soc.ram_encoder_0.current_state\[2\] _1490_ _1502_ _2490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_88_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3498_ _1011_ _1097_ _1098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_25_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5168_ soc.rom_encoder_0.request_data_out\[11\] _2394_ _2437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_56_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4119_ _0954_ _1664_ _1666_ _1667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_83_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5099_ _1404_ _1427_ _2380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_56_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_33_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_70_wb_clk_i clknet_4_12_0_wb_clk_i clknet_leaf_70_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_121_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4470_ soc.spi_video_ram_1.state_counter\[9\] _1975_ _1977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_143_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3421_ _0884_ _1024_ _1025_ soc.cpu.PC.in\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_7_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_98_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3352_ _0945_ _0952_ _0955_ _0875_ _0960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XTAP_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6140_ _0020_ clknet_leaf_1_wb_clk_i soc.video_generator_1.h_count\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_98_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3283_ _0887_ soc.cpu.AReg.data\[1\] _0889_ _0893_ _0894_ _0895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
X_6071_ soc.spi_video_ram_1.write_fifo.fifo_mem\[2\]\[9\] soc.spi_video_ram_1.fifo_in_data\[9\]
+ _3020_ _3030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5022_ _2335_ _1516_ _1529_ soc.ram_encoder_0.request_data_out\[12\] _2336_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_112_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6973_ net53 net50 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5924_ _2949_ _2943_ _2950_ _0570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5855_ _2909_ _0542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_80_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4806_ _0749_ _2176_ _2182_ _2190_ _0212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_21_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5786_ _2846_ _2857_ _2858_ _2849_ _0523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
Xclkbuf_4_15_0_wb_clk_i clknet_0_wb_clk_i clknet_4_15_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_4737_ soc.rom_encoder_0.request_address\[8\] _1650_ _2125_ soc.rom_encoder_0.output_buffer\[5\]
+ _2136_ _2137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_4668_ soc.rom_encoder_0.write_enable _2089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_6407_ _0280_ clknet_leaf_21_wb_clk_i soc.rom_encoder_0.request_address\[12\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3619_ _1216_ _1196_ _1217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_134_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4599_ _2052_ _0142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_88_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6338_ _0213_ clknet_leaf_136_wb_clk_i soc.spi_video_ram_1.buffer_index\[5\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_76_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6269_ _0144_ clknet_leaf_101_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[7\]\[27\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_130_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3970_ soc.ram_encoder_0.output_buffer\[6\] _1520_ _1530_ soc.ram_encoder_0.request_data_out\[2\]
+ _1537_ _1538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_51_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5640_ soc.rom_loader.current_address\[11\] _2767_ _2768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_79_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5571_ soc.spi_video_ram_1.fifo_in_address\[1\] _2705_ _2726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_144_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4522_ soc.spi_video_ram_1.fifo_in_data\[6\] _2007_ _2011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4453_ soc.spi_video_ram_1.state_counter\[3\] _1963_ _1966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_116_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3404_ _0850_ soc.cpu.ALU.x\[8\] _1009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_98_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4384_ _1580_ _1907_ _1908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6123_ _1039_ _2896_ _3052_ _2561_ _0667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_3335_ _0925_ _0935_ _0944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_59_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_58_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3266_ soc.cpu.instruction\[5\] _0879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6054_ _3021_ _0629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5005_ _2322_ soc.rom_encoder_0.request_address\[11\] _2271_ _2323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3197_ _0758_ _0810_ _0811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_82_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_54_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1719 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1708 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5907_ net79 _2936_ _2861_ _2939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_22_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5838_ _2898_ soc.hack_clk_strobe _2893_ _2899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_22_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5769_ soc.cpu.DMuxJMP.sel\[2\] _1669_ _2840_ _2844_ _0846_ _2845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
XFILLER_30_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_89_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_141_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3120_ _0736_ _0008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_95_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6810_ _0652_ clknet_leaf_106_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[2\]\[23\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_24_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3953_ soc.ram_encoder_0.output_buffer\[6\] _1522_ _1525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_91_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6741_ _0583_ clknet_leaf_73_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[0\]\[12\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_51_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6672_ _0514_ clknet_leaf_105_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[6\]\[24\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3884_ soc.video_generator_1.h_count\[2\] _1281_ soc.video_generator_1.h_count\[3\]
+ _1465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_137_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5623_ soc.rom_loader.current_address\[5\] _2755_ _2757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_52_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5554_ soc.spi_video_ram_1.fifo_in_data\[9\] _2708_ _2717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5485_ soc.ram_encoder_0.request_write _2490_ _2530_ _2671_ _2672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_4505_ _1984_ _2000_ _2001_ _0099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_117_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_104_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4436_ soc.spi_video_ram_1.write_fifo.read_pointer\[1\] _1952_ _1954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_116_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4367_ soc.spi_video_ram_1.write_fifo.fifo_mem\[7\]\[14\] _1892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3318_ _0887_ _0927_ _0928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_58_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6106_ soc.spi_video_ram_1.write_fifo.fifo_mem\[2\]\[26\] soc.spi_video_ram_1.fifo_in_address\[10\]
+ _3019_ _3048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xclkbuf_leaf_127_wb_clk_i clknet_4_3_0_wb_clk_i clknet_leaf_127_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_86_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4298_ soc.spi_video_ram_1.write_fifo.fifo_mem\[0\]\[11\] soc.spi_video_ram_1.write_fifo.fifo_mem\[1\]\[11\]
+ soc.spi_video_ram_1.write_fifo.fifo_mem\[2\]\[11\] soc.spi_video_ram_1.write_fifo.fifo_mem\[3\]\[11\]
+ _1584_ _1710_ _1826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3249_ soc.cpu.AReg.data\[1\] _0861_ _0862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_55_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6037_ _3011_ _0622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_23_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_10_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_92_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_72_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5270_ _2514_ _2504_ _2515_ _0351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_114_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4221_ soc.spi_video_ram_1.write_fifo.fifo_mem\[4\]\[6\] soc.spi_video_ram_1.write_fifo.fifo_mem\[5\]\[6\]
+ _1600_ _1754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_68_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4152_ _1581_ _1687_ _1690_ _0685_ _1691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_4083_ _1493_ _1490_ _1504_ _1637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_68_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3103_ _0710_ _0714_ _0719_ _0722_ _0723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_37_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4985_ soc.cpu.PC.REG.data\[6\] soc.rom_loader.current_address\[6\] _2292_ _2308_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_63_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3936_ _0674_ _1492_ _1508_ _1509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
X_6724_ _0566_ net90 net80 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_109_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3867_ _1413_ _1451_ _1452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_20_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6655_ _0497_ clknet_leaf_126_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[6\]\[7\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5606_ _2089_ soc.rom_loader.was_loading _2745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_6586_ net23 clknet_leaf_94_wb_clk_i soc.rom_encoder_0.data_out\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3798_ soc.spi_video_ram_1.output_buffer\[19\] soc.spi_video_ram_1.output_buffer\[16\]
+ soc.spi_video_ram_1.output_buffer\[17\] soc.spi_video_ram_1.output_buffer\[18\]
+ _0757_ _0758_ _1389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_5537_ _2704_ _2708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_133_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_105_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5468_ _2471_ _2658_ _0406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_120_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5399_ _2602_ _2604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_87_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4419_ soc.spi_video_ram_1.write_fifo.fifo_mem\[0\]\[19\] soc.spi_video_ram_1.write_fifo.fifo_mem\[1\]\[19\]
+ soc.spi_video_ram_1.write_fifo.fifo_mem\[2\]\[19\] soc.spi_video_ram_1.write_fifo.fifo_mem\[3\]\[19\]
+ _1594_ _1588_ _1939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_115_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_143_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2025 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2014 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2003 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2058 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2036 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2047 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_95_wb_clk_i clknet_4_11_0_wb_clk_i clknet_leaf_95_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_15_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2069 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_24_wb_clk_i clknet_4_4_0_wb_clk_i clknet_leaf_24_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_42_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput19 la_data_in[10] net19 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_11_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xcaravel_hack_soc_221 wbs_dat_o[28] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xcaravel_hack_soc_210 wbs_dat_o[17] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_6_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_34_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1891 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4770_ _1671_ _2161_ _2162_ _0204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_60_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3721_ _1261_ _1307_ _1319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3652_ _1188_ _1200_ _1250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6440_ _0313_ clknet_leaf_100_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[3\]\[26\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_127_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_115_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6371_ _0244_ clknet_leaf_21_wb_clk_i soc.rom_encoder_0.input_buffer\[5\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_61_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3583_ soc.video_generator_1.v_count\[4\] _1129_ _1181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5322_ soc.ram_encoder_0.request_data_out\[5\] _2545_ _2554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_115_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5253_ soc.ram_encoder_0.toggled_sram_sck _2488_ _2503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_69_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5184_ soc.rom_encoder_0.request_data_out\[15\] _2394_ _2449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4204_ _1711_ _1737_ _1702_ _1738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4135_ soc.ram_encoder_0.output_buffer\[4\] _1509_ _1678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4066_ _1581_ _1614_ _1621_ _1609_ _1622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_36_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4968_ soc.cpu.PC.REG.data\[1\] soc.rom_loader.current_address\[1\] _2293_ _2296_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_51_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3919_ _1488_ _1491_ _1492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_6707_ _0549_ clknet_leaf_53_wb_clk_i soc.ram_encoder_0.address\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4899_ soc.rom_encoder_0.input_buffer\[0\] _2243_ _2250_ _2253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_125_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6638_ _0480_ net89 soc.cpu.ALU.x\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_20_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6569_ _0442_ clknet_leaf_86_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[5\]\[17\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_leaf_142_wb_clk_i clknet_4_0_0_wb_clk_i clknet_leaf_142_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_106_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_11_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_124_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5940_ soc.spi_video_ram_1.write_fifo.fifo_mem\[0\]\[6\] soc.spi_video_ram_1.fifo_in_data\[6\]
+ _2953_ _2960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_53_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5871_ _0745_ _2903_ _2917_ _0550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4822_ _2198_ _0220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_15_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4753_ soc.rom_encoder_0.request_data_out\[5\] _1481_ _2149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_30_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3704_ _1280_ _1301_ _1288_ _1302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_30_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6423_ _0296_ clknet_leaf_81_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[3\]\[9\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4684_ _2100_ _2101_ _0178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3635_ _1175_ _1231_ _1233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_143_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6354_ _0008_ clknet_leaf_133_wb_clk_i soc.spi_video_ram_1.fifo_read_request vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3566_ soc.video_generator_1.v_count\[2\] soc.video_generator_1.v_count\[1\] _1164_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_5305_ _2537_ _2542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_102_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3497_ _0907_ soc.cpu.AReg.data\[13\] _1012_ soc.ram_data_out\[13\] _1097_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6285_ _0160_ clknet_leaf_89_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[4\]\[14\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_130_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5236_ _2487_ soc.ram_encoder_0.input_bits_left\[3\] soc.ram_encoder_0.input_bits_left\[4\]
+ _2488_ _2489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XFILLER_102_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5167_ _0690_ _2436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_97_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4118_ _0923_ _1665_ _1666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_56_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5098_ _2379_ _0315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_29_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4049_ _1592_ _1599_ _1604_ _1605_ _1606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_37_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_65_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_80_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_109_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_48_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_43_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3420_ _0845_ _0926_ soc.cpu.AReg.data\[8\] _0881_ _1025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_3351_ _0884_ _0958_ _0959_ soc.cpu.PC.in\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_48_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3282_ soc.cpu.ALU.zy _0894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XTAP_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6070_ _3029_ _0637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5021_ _1488_ _2334_ _2335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_79_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6972_ net49 net48 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_80_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5923_ soc.gpio_i_stored\[3\] _2943_ _2531_ _2950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_94_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5854_ soc.ram_encoder_0.address\[5\] soc.cpu.AReg.data\[5\] _2903_ _2909_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_21_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4805_ _0720_ _0754_ _2176_ _2189_ _2190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_21_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5785_ soc.cpu.PC.in\[3\] _2851_ _2858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_119_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_108_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4736_ soc.rom_encoder_0.request_data_out\[1\] _1481_ _2136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_4667_ _2088_ _0174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6406_ _0279_ clknet_leaf_21_wb_clk_i soc.rom_encoder_0.request_address\[11\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3618_ soc.display_clks_before_active\[0\] _1216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_115_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4598_ soc.spi_video_ram_1.fifo_in_address\[9\] soc.spi_video_ram_1.write_fifo.fifo_mem\[7\]\[25\]
+ _2037_ _2052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6337_ _0212_ clknet_leaf_112_wb_clk_i soc.spi_video_ram_1.buffer_index\[4\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_1_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3549_ _1141_ _1145_ _1146_ _1147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_131_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6268_ _0143_ clknet_leaf_103_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[7\]\[26\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_103_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5219_ _1403_ _1409_ _2476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6199_ _0079_ clknet_leaf_114_wb_clk_i _0002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_28_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_29_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_63_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5570_ _1597_ _2707_ _2725_ _0441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_102_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4521_ _0009_ _0970_ _2010_ _0106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_8_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4452_ soc.spi_video_ram_1.state_counter\[3\] _1963_ _1965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_3403_ _1000_ _1006_ _1007_ _1008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
X_4383_ _1906_ _1907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_113_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6122_ _1024_ _2896_ _3052_ _2559_ _0666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_3334_ _0884_ _0942_ _0943_ soc.cpu.PC.in\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3265_ soc.cpu.ALU.no _0876_ _0877_ _0878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_2
X_6053_ soc.spi_video_ram_1.write_fifo.fifo_mem\[2\]\[0\] soc.spi_video_ram_1.fifo_in_data\[0\]
+ _3020_ _3021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5004_ soc.cpu.PC.REG.data\[11\] soc.rom_loader.current_address\[11\] _2292_ _2322_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_67_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_66_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3196_ _0759_ _0810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_1709 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5906_ _0902_ _2936_ _2938_ _0564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_34_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5837_ net85 _2898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5768_ _2841_ _2842_ _2843_ _1669_ _2844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_10_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4719_ _1482_ _2123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_5_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5699_ soc.spi_video_ram_1.write_fifo.fifo_mem\[6\]\[3\] soc.spi_video_ram_1.fifo_in_data\[3\]
+ _2799_ _2803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xclkbuf_leaf_49_wb_clk_i clknet_4_6_0_wb_clk_i clknet_leaf_49_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_100_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_130_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_72_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_26_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_107_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6740_ _0582_ clknet_leaf_92_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[0\]\[11\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_23_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3952_ soc.ram_encoder_0.request_address\[5\] _1514_ _1520_ soc.ram_encoder_0.output_buffer\[2\]
+ _1524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_16_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6671_ _0513_ clknet_leaf_104_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[6\]\[23\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_31_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3883_ soc.video_generator_1.h_count\[3\] soc.video_generator_1.h_count\[2\] _1281_
+ _1464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_5622_ soc.rom_loader.current_address\[5\] _2755_ _2756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_31_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5553_ _1787_ _2707_ _2716_ _0433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_129_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4504_ _1128_ _1998_ _2001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5484_ _1512_ _2670_ _2671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4435_ soc.spi_video_ram_1.write_fifo.read_pointer\[1\] _1952_ _1953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4366_ _1600_ soc.spi_video_ram_1.write_fifo.fifo_mem\[4\]\[14\] _1890_ _1891_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_141_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3317_ soc.ram_data_out\[3\] _0869_ _0927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_86_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_86_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6105_ _3047_ _0654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_112_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4297_ _1575_ _1611_ _1825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3248_ soc.cpu.AReg.data\[3\] soc.cpu.AReg.data\[2\] _0861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6036_ soc.spi_video_ram_1.fifo_in_address\[6\] soc.spi_video_ram_1.write_fifo.fifo_mem\[1\]\[22\]
+ _2999_ _3011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_132_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3179_ _0762_ _0786_ _0792_ _0780_ _0793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_26_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_14_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_35 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_131_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_65_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_61_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_14_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_13_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_139_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4220_ _1592_ _1750_ _1752_ _1605_ _1753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_123_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4151_ _1605_ _1689_ _1690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4082_ _1497_ soc.ram_encoder_0.output_bits_left\[4\] _1636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_110_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3102_ _0720_ _0721_ _0722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_110_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4984_ _2307_ _0273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_23_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3935_ _1493_ _1495_ _1496_ _1507_ _1508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
X_6723_ _0565_ net90 net79 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6654_ _0496_ clknet_leaf_123_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[6\]\[6\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5605_ soc.rom_loader.current_address\[0\] _0473_ _2744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_3866_ soc.rom_encoder_0.output_buffer\[19\] _1417_ _1442_ soc.rom_encoder_0.request_data_out\[15\]
+ _1451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_31_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6585_ net22 clknet_leaf_94_wb_clk_i soc.rom_encoder_0.data_out\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3797_ _1381_ _1383_ _1387_ _1388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_106_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5536_ _2704_ _2707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_117_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5467_ soc.ram_data_out\[14\] _2604_ _2657_ _2658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4418_ _1578_ _1937_ _1938_ _0075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_114_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5398_ _2602_ _2603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_28_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_143_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_87_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4349_ _0729_ _1181_ _1874_ _1875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_143_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6019_ _1860_ _2988_ _3002_ _0613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_2015 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2004 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2059 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2037 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2048 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2026 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_139_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_64_wb_clk_i clknet_4_12_0_wb_clk_i clknet_leaf_64_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_10_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_6_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xcaravel_hack_soc_222 wbs_dat_o[29] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_10_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xcaravel_hack_soc_200 wbs_dat_o[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xcaravel_hack_soc_211 wbs_dat_o[18] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_123_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_92_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1870 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1892 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1881 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3720_ _1236_ _1317_ _1318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_9_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3651_ soc.video_generator_1.h_count\[9\] _1134_ _1249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_6370_ _0243_ clknet_leaf_18_wb_clk_i soc.rom_encoder_0.input_buffer\[4\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3582_ _1157_ _1161_ _1178_ _1179_ _1180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_138_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5321_ soc.ram_encoder_0.data_out\[5\] _2553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_54_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5252_ soc.ram_encoder_0.input_buffer\[0\] _2502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_142_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5183_ _2436_ _2448_ _0331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4203_ soc.spi_video_ram_1.write_fifo.fifo_mem\[2\]\[5\] soc.spi_video_ram_1.write_fifo.fifo_mem\[3\]\[5\]
+ _1600_ _1737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4134_ soc.ram_encoder_0.request_address\[3\] _1514_ _1677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_111_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_56_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4065_ _1592_ _1617_ _1620_ _1605_ _1621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_3_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4967_ _2295_ _0268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3918_ _1489_ _1490_ _1491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_6706_ _0548_ clknet_leaf_70_wb_clk_i soc.ram_encoder_0.address\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4898_ soc.rom_encoder_0.input_buffer\[4\] _2252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6637_ _0479_ net89 soc.cpu.ALU.x\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3849_ _1412_ _1434_ _1435_ _1436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_6568_ _0441_ clknet_leaf_83_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[5\]\[16\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5519_ _2691_ _2694_ _2695_ _0420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_4_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6499_ _0372_ clknet_leaf_49_wb_clk_i soc.ram_encoder_0.request_data_out\[12\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_105_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_111_wb_clk_i clknet_4_8_0_wb_clk_i clknet_leaf_111_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_59_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_31_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_11_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_111_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_120_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5870_ soc.ram_encoder_0.address\[13\] _2903_ _2917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_74_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4821_ soc.spi_video_ram_1.fifo_in_address\[5\] soc.cpu.AReg.data\[5\] _2018_ _2198_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_2390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4752_ _2122_ _2147_ _2148_ _0200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_105_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4683_ soc.spi_video_ram_1.state_sram_clk_counter\[2\] _2098_ _2096_ _2101_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3703_ soc.video_generator_1.h_count\[3\] _1196_ _1269_ _1301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_88_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3634_ _1175_ _1231_ _1232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_6422_ _0295_ clknet_leaf_114_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[3\]\[8\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_134_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6353_ _0227_ clknet_leaf_79_wb_clk_i soc.spi_video_ram_1.fifo_in_address\[12\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_3565_ _1125_ _1162_ _1128_ _1148_ _1163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_115_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5304_ soc.ram_encoder_0.data_out\[0\] _2541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_103_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3496_ _0923_ _1095_ _1096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_6284_ _0159_ clknet_leaf_87_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[4\]\[13\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5235_ soc.ram_encoder_0.current_state\[2\] _1496_ _2488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_103_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5166_ _2400_ _2435_ _0327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_29_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4117_ _0904_ soc.cpu.ALU.x\[15\] _1665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_57_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5097_ soc.spi_video_ram_1.write_fifo.fifo_mem\[3\]\[28\] soc.spi_video_ram_1.fifo_in_address\[12\]
+ _2216_ _2379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4048_ _1579_ _1605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_44_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_140_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_5999_ soc.spi_video_ram_1.fifo_in_data\[4\] soc.spi_video_ram_1.write_fifo.fifo_mem\[1\]\[4\]
+ _2986_ _2992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_40_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_16_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3350_ _0846_ soc.cpu.instruction\[4\] soc.cpu.AReg.data\[4\] _0881_ _0959_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_98_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5020_ _1493_ soc.ram_encoder_0.current_state\[1\] _2334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_112_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3281_ _0890_ _0868_ _0891_ _0892_ _0869_ _0893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XTAP_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6971_ net49 net47 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_65_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5922_ net17 _2949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_94_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5853_ _2908_ _0541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_80_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_22_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_142_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5784_ soc.cpu.PC.REG.data\[3\] _2856_ _2857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_10_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4804_ _0720_ _1383_ _2189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_22_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4735_ _2122_ _2134_ _2135_ _0196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_107_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4666_ soc.spi_video_ram_1.write_fifo.fifo_mem\[4\]\[28\] soc.spi_video_ram_1.fifo_in_address\[12\]
+ _2057_ _2088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_135_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6405_ _0278_ clknet_leaf_29_wb_clk_i soc.rom_encoder_0.request_address\[10\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4597_ _2051_ _0141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3617_ soc.video_generator_1.h_count\[3\] _1196_ _1215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6336_ _0211_ clknet_leaf_136_wb_clk_i soc.spi_video_ram_1.buffer_index\[3\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3548_ soc.boot_loading_offset\[1\] _1144_ _1146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_89_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3479_ _1005_ _1008_ _1079_ _1080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_76_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6267_ _0142_ clknet_leaf_111_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[7\]\[25\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5218_ _2380_ _2474_ _2475_ _2471_ _0339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_6198_ _0078_ clknet_leaf_133_wb_clk_i _0001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_97_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5149_ _0990_ _2392_ _2422_ _2423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_57_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_31_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4520_ soc.spi_video_ram_1.fifo_in_data\[5\] _2007_ _2010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_117_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4451_ _1961_ _1963_ _1964_ _0082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_144_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3402_ _0986_ _0999_ _1007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6121_ _1002_ _2897_ _3052_ _2557_ _0665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XTAP_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4382_ soc.spi_video_ram_1.write_fifo.fifo_mem\[4\]\[23\] soc.spi_video_ram_1.write_fifo.fifo_mem\[5\]\[23\]
+ soc.spi_video_ram_1.write_fifo.fifo_mem\[6\]\[23\] soc.spi_video_ram_1.write_fifo.fifo_mem\[7\]\[23\]
+ _1582_ _0001_ _1906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_112_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3333_ _0845_ soc.cpu.instruction\[3\] soc.cpu.AReg.data\[3\] _0881_ _0943_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai22_1
XTAP_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3264_ _0852_ _0874_ _0877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6052_ _3019_ _3020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_5003_ _2272_ _2320_ _2321_ _0278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_78_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3195_ soc.spi_video_ram_1.output_buffer\[8\] soc.spi_video_ram_1.output_buffer\[9\]
+ _0783_ _0809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_22_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5905_ net78 _2936_ _2861_ _2938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_81_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5836_ _2896_ _2897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_50_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5767_ _1069_ _1108_ _2838_ _2843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_50_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4718_ _1670_ _2122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_5698_ _2802_ _0492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_108_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4649_ _2079_ _0165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_89_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_131_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6319_ _0194_ clknet_leaf_25_wb_clk_i soc.rom_encoder_0.output_buffer\[6\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_1_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_103_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_89_wb_clk_i clknet_4_11_0_wb_clk_i clknet_leaf_89_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
Xclkbuf_leaf_18_wb_clk_i clknet_4_4_0_wb_clk_i clknet_leaf_18_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_58_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_91_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_73_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_99_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3951_ _1510_ _1521_ _1523_ _0024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_50_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3882_ soc.video_generator_1.h_count\[2\] _1281_ _1463_ _0015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_32_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6670_ _0512_ clknet_leaf_97_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[6\]\[22\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5621_ _2746_ _2754_ _2755_ _0461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_84_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5552_ soc.spi_video_ram_1.fifo_in_data\[8\] _2708_ _2716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4503_ soc.video_generator_1.v_count\[8\] _1999_ _2000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5483_ _2601_ _2668_ _2669_ _2670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_105_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4434_ _1461_ _1951_ _1952_ _0077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_113_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4365_ _1593_ _1889_ _1890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_140_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3316_ _0853_ _0926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_59_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6104_ soc.spi_video_ram_1.write_fifo.fifo_mem\[2\]\[25\] soc.spi_video_ram_1.fifo_in_address\[9\]
+ _3019_ _3047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_100_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6035_ _3010_ _0621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4296_ _1811_ _1823_ _1824_ _0067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_101_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3247_ _0856_ _0857_ _0858_ _0859_ _0860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_73_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3178_ _0775_ _0787_ _0791_ _0762_ _0792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_27_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_26_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xclkbuf_leaf_136_wb_clk_i clknet_4_2_0_wb_clk_i clknet_leaf_136_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_22_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5819_ _2846_ _2882_ _2883_ _0531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_109_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6799_ _0641_ clknet_leaf_74_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[2\]\[12\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_136_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_61_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_41_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4150_ _1688_ _1689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_95_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3101_ soc.spi_video_ram_1.state_sram_clk_counter\[2\] _0713_ _0721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4081_ _1634_ _1635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_96_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_64_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4983_ _2306_ soc.rom_encoder_0.request_address\[5\] _2287_ _2307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_51_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3934_ soc.ram_encoder_0.toggled_sram_sck _1506_ _1507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_108_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6722_ _0564_ net88 net78 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_51_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6653_ _0495_ clknet_leaf_124_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[6\]\[5\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_32_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3865_ _1432_ _1449_ _1450_ _0676_ _0011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_5604_ _1403_ _0691_ _0456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_118_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6584_ net21 clknet_leaf_27_wb_clk_i soc.rom_encoder_0.data_out\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3796_ _1384_ _1386_ _1387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_20_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5535_ _2706_ _0425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_11_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5466_ _2526_ _2606_ _2602_ _2656_ _2657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_4417_ soc.spi_video_ram_1.output_buffer\[5\] _1611_ _1938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5397_ _1489_ soc.ram_encoder_0.current_state\[1\] _2601_ _2602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_99_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4348_ _0686_ _1859_ _1873_ _1850_ _1874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4279_ _1802_ _1808_ _1809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_47_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6018_ soc.spi_video_ram_1.fifo_in_data\[13\] _2986_ _3002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_2016 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2005 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2038 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2049 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2027 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xcaravel_hack_soc_201 wbs_dat_o[8] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_108_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xcaravel_hack_soc_223 wbs_dat_o[30] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xcaravel_hack_soc_212 wbs_dat_o[19] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_124_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xclkbuf_leaf_33_wb_clk_i clknet_4_5_0_wb_clk_i clknet_leaf_33_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_123_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1860 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1893 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1882 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1871 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3650_ _1176_ _1186_ _1246_ _1248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_3581_ soc.boot_loading_offset\[3\] _1177_ _1179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_115_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5320_ _2551_ _2542_ _2552_ _0364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_6_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5251_ _2498_ _2500_ _2501_ _0346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_102_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4202_ _1595_ soc.spi_video_ram_1.write_fifo.fifo_mem\[0\]\[5\] _1735_ _1736_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_123_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5182_ soc.cpu.instruction\[14\] _2393_ _2447_ _2448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_110_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4133_ _1676_ _0052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_69_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4064_ _1601_ soc.spi_video_ram_1.write_fifo.fifo_mem\[6\]\[18\] _1619_ _1588_ _1620_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_25_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6705_ _0547_ clknet_leaf_70_wb_clk_i soc.ram_encoder_0.address\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4966_ _2294_ soc.rom_encoder_0.request_address\[0\] _2287_ _2295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3917_ soc.ram_encoder_0.current_state\[1\] _1490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_4897_ _2249_ _2242_ _2251_ _0242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_6636_ _0478_ net89 soc.cpu.ALU.x\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3848_ _1426_ _1419_ _1435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_22_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6567_ _0440_ clknet_leaf_72_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[5\]\[15\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3779_ _0836_ _1370_ _1364_ _1371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_118_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5518_ soc.hack_clock_0.counter\[2\] _2693_ _2695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xclkbuf_4_1_0_wb_clk_i clknet_0_wb_clk_i clknet_4_1_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_118_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6498_ _0371_ clknet_leaf_46_wb_clk_i soc.ram_encoder_0.request_data_out\[11\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5449_ soc.ram_encoder_0.request_data_out\[10\] _2605_ _2644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_78_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4820_ _2197_ _0219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_61_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4751_ soc.rom_encoder_0.output_buffer\[12\] _2138_ _2148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_30_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4682_ soc.spi_video_ram_1.state_sram_clk_counter\[2\] _2098_ _2100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_3702_ _1278_ _1296_ _1299_ _1286_ _1300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_30_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3633_ _1195_ _1198_ _1231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_6421_ _0294_ clknet_leaf_127_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[3\]\[7\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_115_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6352_ _0226_ clknet_leaf_76_wb_clk_i soc.spi_video_ram_1.fifo_in_address\[11\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_3564_ soc.video_generator_1.v_count\[3\] _1162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_115_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5303_ _2538_ _2539_ _2540_ _0359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3495_ _0904_ soc.cpu.ALU.x\[13\] _1095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6283_ _0158_ clknet_leaf_93_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[4\]\[12\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_143_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_142_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5234_ soc.ram_encoder_0.input_bits_left\[2\] _2487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_102_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5165_ _0923_ _2393_ _2434_ _2435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_111_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4116_ _0926_ _1663_ _1664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_25_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5096_ _2378_ _0314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_83_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_72_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4047_ _1601_ soc.spi_video_ram_1.write_fifo.fifo_mem\[6\]\[16\] _1603_ _1588_ _1604_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_24_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_25_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_80_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_52_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5998_ _2991_ _0603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4949_ _2284_ _0261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_71_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6619_ soc.cpu.PC.in\[2\] net87 soc.cpu.AReg.data\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_4_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_121_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_90_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_16_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_7_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_124_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3280_ soc.gpio_i_stored\[1\] _0855_ _0860_ _0865_ _0892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6970_ net49 net46 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_81_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_54_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5921_ _2947_ _2943_ _2948_ _0569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_47_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5852_ soc.ram_encoder_0.address\[4\] soc.cpu.AReg.data\[4\] _2903_ _2908_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_62_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5783_ soc.cpu.PC.REG.data\[0\] soc.cpu.PC.REG.data\[1\] soc.cpu.PC.REG.data\[2\]
+ _2856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_4803_ _1796_ _2188_ _0211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_21_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4734_ soc.rom_encoder_0.output_buffer\[8\] _1671_ _2135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_30_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4665_ _2087_ _0173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6404_ _0277_ clknet_leaf_20_wb_clk_i soc.rom_encoder_0.request_address\[9\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4596_ soc.spi_video_ram_1.fifo_in_address\[8\] soc.spi_video_ram_1.write_fifo.fifo_mem\[7\]\[24\]
+ _2037_ _2051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3616_ _1208_ _1212_ _1213_ _1214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_6335_ _0210_ clknet_leaf_136_wb_clk_i soc.spi_video_ram_1.buffer_index\[2\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3547_ soc.boot_loading_offset\[1\] _1144_ _1145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_142_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_103_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3478_ _1078_ _1079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6266_ _0141_ clknet_leaf_105_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[7\]\[24\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5217_ _1438_ _2380_ soc.rom_encoder_0.initializing_step\[1\] _2475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_6197_ _0077_ clknet_leaf_133_wb_clk_i _0000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_96_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5148_ _2247_ _2413_ _2414_ _2421_ _2422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_5079_ soc.spi_video_ram_1.write_fifo.fifo_mem\[3\]\[19\] soc.spi_video_ram_1.fifo_in_address\[3\]
+ _2368_ _2370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_72_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_5_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4450_ soc.spi_video_ram_1.state_counter\[1\] soc.spi_video_ram_1.state_counter\[0\]
+ soc.spi_video_ram_1.state_counter\[2\] _1964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3401_ _0983_ _1004_ _1006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_4381_ soc.spi_video_ram_1.write_fifo.fifo_mem\[0\]\[23\] soc.spi_video_ram_1.write_fifo.fifo_mem\[1\]\[23\]
+ soc.spi_video_ram_1.write_fifo.fifo_mem\[2\]\[23\] soc.spi_video_ram_1.write_fifo.fifo_mem\[3\]\[23\]
+ _1755_ _1587_ _1905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_113_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6120_ _0989_ _2897_ _3052_ _2555_ _0664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_3332_ _0922_ _0941_ _0942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_98_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3263_ _0852_ _0874_ _0875_ _0876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6051_ _3018_ _3019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_112_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5002_ soc.rom_encoder_0.request_address\[10\] _2272_ _2321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3194_ _0758_ _0759_ _0808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XTAP_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5904_ _0878_ _2936_ _2937_ _0563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5835_ _2895_ _2896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_22_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5766_ _0990_ _1122_ _2842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_5697_ soc.spi_video_ram_1.write_fifo.fifo_mem\[6\]\[2\] soc.spi_video_ram_1.fifo_in_data\[2\]
+ _2799_ _2802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4717_ _2121_ _0192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_135_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4648_ soc.spi_video_ram_1.write_fifo.fifo_mem\[4\]\[19\] soc.spi_video_ram_1.fifo_in_address\[3\]
+ _2069_ _2079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_30_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4579_ _2042_ _0132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_1_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6318_ _0193_ clknet_leaf_25_wb_clk_i soc.rom_encoder_0.output_buffer\[5\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_104_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6249_ _0124_ clknet_leaf_120_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[7\]\[7\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_18_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_84_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_58_wb_clk_i clknet_4_13_0_wb_clk_i clknet_leaf_58_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_72_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_4_14_0_wb_clk_i clknet_0_wb_clk_i clknet_4_14_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_76_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3950_ soc.ram_encoder_0.output_buffer\[5\] _1522_ _1523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_32_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3881_ soc.video_generator_1.h_count\[2\] _1281_ _1462_ _1463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5620_ soc.rom_loader.current_address\[4\] _2753_ _2755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_77_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5551_ _1767_ _2707_ _2715_ _0432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_117_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4502_ _1984_ _1997_ _1999_ _0098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_144_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5482_ _1517_ _2533_ _2669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_104_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4433_ _0697_ _1949_ _0702_ _1952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_99_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4364_ soc.spi_video_ram_1.write_fifo.fifo_mem\[5\]\[14\] _1889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_98_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3315_ _0923_ _0924_ _0925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6103_ _3046_ _0653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4295_ soc.spi_video_ram_1.output_buffer\[13\] _1612_ _1824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3246_ soc.cpu.AReg.data\[9\] soc.cpu.AReg.data\[8\] _0859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_86_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6034_ soc.spi_video_ram_1.fifo_in_address\[5\] soc.spi_video_ram_1.write_fifo.fifo_mem\[1\]\[21\]
+ _2999_ _3010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3177_ _0775_ _0790_ _0791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_27_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_81_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_35_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5818_ soc.cpu.PC.in\[11\] _2847_ _2861_ _2883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6798_ _0640_ clknet_leaf_90_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[2\]\[11\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_50_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5749_ _2828_ _0517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xclkbuf_leaf_105_wb_clk_i clknet_4_10_0_wb_clk_i clknet_leaf_105_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_123_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_85_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput80 net80 io_out[37] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_3100_ soc.spi_video_ram_1.current_state\[3\] _0720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
X_4080_ _0674_ soc.ram_encoder_0.toggled_sram_sck _1506_ _1515_ _1634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_110_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4982_ soc.cpu.PC.REG.data\[5\] soc.rom_loader.current_address\[5\] _2292_ _2306_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_63_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3933_ _1499_ _1505_ _1506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6721_ _0563_ net91 net77 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_60_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_3_wb_clk_i clknet_4_1_0_wb_clk_i clknet_leaf_3_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_108_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6652_ _0494_ clknet_leaf_12_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[6\]\[4\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_32_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3864_ net66 _1432_ _1450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5603_ _1461_ _2742_ _0473_ _0455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_3795_ _1382_ _1385_ _1386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_6583_ net20 clknet_leaf_143_wb_clk_i soc.rom_encoder_0.data_out\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_118_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5534_ soc.spi_video_ram_1.fifo_in_data\[0\] soc.spi_video_ram_1.write_fifo.fifo_mem\[5\]\[0\]
+ _2705_ _2706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_11_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5465_ soc.ram_encoder_0.request_data_out\[14\] _2605_ _2656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_105_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4416_ _1581_ _1929_ _1936_ _1609_ _1937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_132_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5396_ _1504_ _1499_ _2489_ soc.ram_encoder_0.toggled_sram_sck _2601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_113_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4347_ _0703_ _1865_ _1872_ _1873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_4278_ _1711_ _1803_ _1807_ _1808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_86_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6017_ _3001_ _0612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_67_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3229_ soc.spi_video_ram_1.buffer_index\[4\] _0819_ _0842_ _0752_ _0843_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai22_1
XTAP_2006 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2039 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2028 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2017 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xcaravel_hack_soc_202 wbs_dat_o[9] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_136_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xcaravel_hack_soc_224 wbs_dat_o[31] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xcaravel_hack_soc_213 wbs_dat_o[20] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_10_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_78_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_leaf_73_wb_clk_i clknet_4_15_0_wb_clk_i clknet_leaf_73_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_93_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1861 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1850 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1894 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1872 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3580_ soc.boot_loading_offset\[3\] _1177_ _1178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_142_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5250_ soc.ram_encoder_0.input_bits_left\[4\] _2497_ _2501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_114_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4201_ _1601_ _1734_ _1591_ _1735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_69_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5181_ _2264_ _2395_ _2391_ _2446_ _2447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_110_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4132_ soc.rom_encoder_0.output_buffer\[1\] _1671_ _1672_ soc.rom_encoder_0.request_address\[0\]
+ _1676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_3_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4063_ _1594_ _1618_ _1619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_49_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4965_ soc.cpu.PC.REG.data\[0\] soc.rom_loader.current_address\[0\] _2293_ _2294_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3916_ soc.ram_encoder_0.current_state\[2\] _1489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_6704_ _0546_ clknet_leaf_64_wb_clk_i soc.ram_encoder_0.address\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_138_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4896_ net8 _2243_ _2250_ _2251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_60_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6635_ _0477_ net89 soc.cpu.ALU.x\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3847_ soc.rom_encoder_0.output_bits_left\[4\] _1433_ _1434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_20_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6566_ _0439_ clknet_leaf_85_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[5\]\[14\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3778_ _0808_ _0838_ _0760_ _1370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_20_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5517_ soc.hack_clock_0.counter\[2\] _2693_ _2694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_6497_ _0370_ clknet_leaf_43_wb_clk_i soc.ram_encoder_0.request_data_out\[10\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_105_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5448_ _2615_ _2643_ _0401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5379_ _2588_ _0387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_87_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_120_wb_clk_i clknet_4_9_0_wb_clk_i clknet_leaf_120_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_11_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_124_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4750_ soc.rom_encoder_0.request_address\[11\] _1650_ _2125_ soc.rom_encoder_0.output_buffer\[8\]
+ _2146_ _2147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_61_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4681_ _2098_ _2099_ _0177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3701_ _1297_ _1298_ _1299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6420_ _0293_ clknet_leaf_124_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[3\]\[6\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3632_ _1223_ _1228_ _1229_ _1230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_127_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6351_ _0225_ clknet_leaf_75_wb_clk_i soc.spi_video_ram_1.fifo_in_address\[10\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_115_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5302_ soc.ram_encoder_0.request_write _2538_ _2540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3563_ _1158_ _1159_ _1153_ _1160_ _1161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_143_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_143_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3494_ _1076_ _1094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6282_ _0157_ clknet_leaf_95_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[4\]\[11\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5233_ _2436_ soc.ram_encoder_0.toggled_sram_sck _0343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_103_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5164_ _2256_ _2413_ _2414_ _2433_ _2434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_110_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4115_ _1011_ _1662_ _1663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_84_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5095_ soc.spi_video_ram_1.write_fifo.fifo_mem\[3\]\[27\] soc.spi_video_ram_1.fifo_in_address\[11\]
+ _2368_ _2378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_65_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4046_ _1594_ _1602_ _1603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_37_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_25_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_64_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_80_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5997_ soc.spi_video_ram_1.fifo_in_data\[3\] soc.spi_video_ram_1.write_fifo.fifo_mem\[1\]\[3\]
+ _2986_ _2991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4948_ soc.rom_encoder_0.data_out\[9\] soc.rom_encoder_0.request_data_out\[9\] _2276_
+ _2284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_12_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4879_ _2236_ _2237_ _2238_ _0237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_32_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6618_ soc.cpu.PC.in\[1\] net88 soc.cpu.AReg.data\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_21_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6549_ _0422_ clknet_leaf_36_wb_clk_i soc.hack_clock_0.counter\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_106_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_74_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_112_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_66_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5920_ soc.gpio_i_stored\[2\] _2943_ _2531_ _2948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_81_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_81_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5851_ _2907_ _0540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_22_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5782_ _2846_ _2854_ _2855_ _2849_ _0522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_4802_ _0752_ _2185_ _2188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_21_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4733_ soc.rom_encoder_0.request_address\[7\] _1650_ _2125_ soc.rom_encoder_0.output_buffer\[4\]
+ _2133_ _2134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_6403_ _0276_ clknet_leaf_20_wb_clk_i soc.rom_encoder_0.request_address\[8\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4664_ soc.spi_video_ram_1.write_fifo.fifo_mem\[4\]\[27\] soc.spi_video_ram_1.fifo_in_address\[11\]
+ _2057_ _2087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4595_ _2050_ _0140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3615_ _1166_ _1169_ _1158_ _1213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_6334_ _0209_ clknet_leaf_112_wb_clk_i soc.spi_video_ram_1.buffer_index\[1\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3546_ _1142_ soc.video_generator_1.v_count\[1\] _1143_ _1144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_142_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6265_ _0140_ clknet_leaf_104_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[7\]\[23\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_89_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3477_ _1046_ _1048_ _1077_ _1078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_5216_ _2472_ _2473_ _2474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_88_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6196_ _0076_ clknet_leaf_115_wb_clk_i soc.spi_video_ram_1.output_buffer\[4\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_130_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5147_ soc.rom_encoder_0.request_data_out\[6\] _2395_ _2421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_56_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5078_ _2369_ _0305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4029_ _0001_ _1586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_38_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3400_ _0945_ _0981_ _1004_ _1005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_4380_ _1702_ _1900_ _1903_ _1904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3331_ _0875_ _0938_ _0940_ _0941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_124_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3262_ soc.cpu.ALU.f _0875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_2
XTAP_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6050_ soc.spi_video_ram_1.write_fifo.write_pointer\[2\] _2703_ _0698_ _3018_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_112_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5001_ _2293_ soc.rom_loader.current_address\[10\] _2319_ _2320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_66_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3193_ _0720_ soc.spi_video_ram_1.buffer_index\[5\] _0807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_38_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5903_ net77 _2936_ _2861_ _2937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_81_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_81_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5834_ _0744_ _2894_ _2895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_50_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5765_ soc.cpu.DMuxJMP.sel\[1\] _2841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5696_ _2801_ _0491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4716_ net12 soc.spi_video_ram_1.read_value\[3\] _2117_ _2121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4647_ _2078_ _0164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_144_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4578_ soc.spi_video_ram_1.fifo_in_data\[15\] soc.spi_video_ram_1.write_fifo.fifo_mem\[7\]\[15\]
+ _2037_ _2042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6317_ _0192_ clknet_leaf_145_wb_clk_i soc.spi_video_ram_1.read_value\[3\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_1_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3529_ soc.video_generator_1.v_count\[5\] _1127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_6248_ _0123_ clknet_leaf_122_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[7\]\[6\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6179_ _0059_ clknet_leaf_134_wb_clk_i soc.spi_video_ram_1.output_buffer\[21\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_58_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_45_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_98_wb_clk_i clknet_4_11_0_wb_clk_i clknet_leaf_98_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_38_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_27_wb_clk_i clknet_4_5_0_wb_clk_i clknet_leaf_27_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_40_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_96_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3880_ _1460_ _1462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5550_ soc.spi_video_ram_1.fifo_in_data\[7\] _2708_ _2715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_144_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_129_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5481_ _2334_ _1495_ _2667_ _2668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_8_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4501_ _1168_ _1998_ _1999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4432_ soc.spi_video_ram_1.write_fifo.read_pointer\[0\] _1950_ _1951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_126_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4363_ _1885_ _1887_ _1888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_99_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3314_ _0904_ soc.cpu.ALU.x\[3\] _0924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4294_ _0729_ _1813_ _1816_ _1609_ _1822_ _1823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_6102_ soc.spi_video_ram_1.write_fifo.fifo_mem\[2\]\[24\] soc.spi_video_ram_1.fifo_in_address\[8\]
+ _3019_ _3046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_141_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_98_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3245_ soc.cpu.AReg.data\[14\] soc.cpu.AReg.data\[13\] _0858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_86_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6033_ _3009_ _0620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_6_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3176_ _0771_ _0788_ _0789_ _0757_ _0790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_94_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_82_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_22_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5817_ soc.cpu.PC.REG.data\[11\] _2881_ _2882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_6797_ _0639_ clknet_leaf_91_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[2\]\[10\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_50_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5748_ soc.spi_video_ram_1.write_fifo.fifo_mem\[6\]\[27\] soc.spi_video_ram_1.fifo_in_address\[11\]
+ _2798_ _2828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_135_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5679_ _1058_ _2779_ _2791_ _0484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_68_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_145_wb_clk_i clknet_4_0_0_wb_clk_i clknet_leaf_145_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_104_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xoutput70 net70 io_out[22] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_123_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_110_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput81 net81 io_out[8] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_110_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4981_ _2305_ _0272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_45_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3932_ soc.ram_encoder_0.request_write _1501_ _1504_ _1505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6720_ _0562_ clknet_leaf_8_wb_clk_i soc.hack_wait_clocks\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6651_ _0493_ clknet_leaf_15_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[6\]\[3\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3863_ soc.rom_encoder_0.output_buffer\[18\] _1436_ _1448_ _1441_ _1449_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_5602_ _2743_ _0473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6582_ _0455_ clknet_leaf_6_wb_clk_i soc.rom_loader.writing vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5533_ _2704_ _2705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
X_3794_ _0759_ _0764_ _0752_ _1385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_117_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5464_ _2471_ _2655_ _0405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5395_ _1461_ _2594_ _2599_ _2600_ _0391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_4415_ _1592_ _1932_ _1935_ _1702_ _1936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_113_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_28_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4346_ _1591_ _1868_ _1871_ _1579_ _1872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_101_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_100_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_86_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4277_ _1580_ _1806_ _1807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6016_ soc.spi_video_ram_1.fifo_in_data\[12\] soc.spi_video_ram_1.write_fifo.fifo_mem\[1\]\[12\]
+ _2999_ _3001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3228_ _0832_ _0841_ _0842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_27_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2007 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3159_ _0757_ soc.spi_video_ram_1.output_buffer\[6\] _0772_ soc.spi_video_ram_1.output_buffer\[7\]
+ _0773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_36_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2029 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2018 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xcaravel_hack_soc_214 wbs_dat_o[21] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xcaravel_hack_soc_203 wbs_dat_o[10] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xcaravel_hack_soc_225 io_oeb[26] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_136_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_77_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_42_wb_clk_i clknet_4_7_0_wb_clk_i clknet_leaf_42_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_34_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1851 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1840 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1884 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1873 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1862 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1895 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4200_ soc.spi_video_ram_1.write_fifo.fifo_mem\[1\]\[5\] _1734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_111_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5180_ soc.rom_encoder_0.request_data_out\[14\] _2394_ _2446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_96_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4131_ _1675_ _0051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_68_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4062_ soc.spi_video_ram_1.write_fifo.fifo_mem\[7\]\[18\] _1618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_92_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4964_ _2292_ _2293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_52_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3915_ soc.ram_encoder_0.current_state\[0\] _1488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
X_6703_ _0545_ clknet_leaf_65_wb_clk_i soc.ram_encoder_0.address\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_32_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4895_ _0675_ _2250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_6634_ _0476_ net89 soc.cpu.ALU.x\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3846_ soc.rom_encoder_0.output_bits_left\[2\] _1415_ _1433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6565_ _0438_ clknet_leaf_87_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[5\]\[13\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3777_ _0776_ soc.spi_video_ram_1.output_buffer\[1\] _0811_ _1369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_6496_ _0369_ clknet_leaf_43_wb_clk_i soc.ram_encoder_0.request_data_out\[9\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5516_ _2691_ _2692_ _2693_ _0419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_118_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5447_ soc.ram_data_out\[9\] _2603_ _2642_ _2643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_121_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5378_ soc.ram_encoder_0.address\[11\] soc.ram_encoder_0.request_address\[11\] _2581_
+ _2588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_87_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4329_ soc.spi_video_ram_1.write_fifo.fifo_mem\[0\]\[25\] soc.spi_video_ram_1.write_fifo.fifo_mem\[1\]\[25\]
+ soc.spi_video_ram_1.write_fifo.fifo_mem\[2\]\[25\] soc.spi_video_ram_1.write_fifo.fifo_mem\[3\]\[25\]
+ _1755_ _1590_ _1855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_101_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_34_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1692 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3700_ _1216_ _1218_ _1219_ _1298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4680_ soc.spi_video_ram_1.state_sram_clk_counter\[1\] _2095_ _2096_ _2099_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3631_ _1225_ _1227_ _1229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6350_ _0224_ clknet_leaf_77_wb_clk_i soc.spi_video_ram_1.fifo_in_address\[9\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_3562_ soc.boot_loading_offset\[1\] _1144_ _1160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_115_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5301_ soc.synch_hack_writeM _0869_ _2539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_52_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3493_ _0883_ _1092_ _1093_ soc.cpu.PC.in\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_6281_ _0156_ clknet_leaf_90_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[4\]\[10\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_130_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5232_ soc.rom_encoder_0.initializing_step\[4\] _2484_ _2486_ _2471_ _0342_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_5163_ soc.rom_encoder_0.request_data_out\[10\] _2394_ _2433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_96_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4114_ _0907_ soc.cpu.AReg.data\[15\] _1012_ soc.ram_data_out\[15\] _1662_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_111_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5094_ _2377_ _0313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4045_ soc.spi_video_ram_1.write_fifo.fifo_mem\[7\]\[16\] _1602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_17_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_37_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_80_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5996_ _2990_ _0602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_40_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4947_ _2283_ _0260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_33_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4878_ soc.rom_encoder_0.input_bits_left\[2\] _2232_ soc.rom_encoder_0.input_bits_left\[3\]
+ _2238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_137_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6617_ soc.cpu.PC.in\[0\] net91 soc.cpu.AReg.data\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_3829_ soc.rom_encoder_0.output_bits_left\[2\] _1414_ _1415_ _1416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_20_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6548_ _0421_ clknet_leaf_36_wb_clk_i soc.hack_clock_0.counter\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6479_ _0352_ clknet_leaf_60_wb_clk_i soc.ram_encoder_0.input_buffer\[5\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_133_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_31_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_94_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5850_ soc.ram_encoder_0.address\[3\] soc.cpu.AReg.data\[3\] _2903_ _2907_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_62_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5781_ soc.cpu.PC.in\[2\] _2851_ _2855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4801_ _2182_ _2185_ _2187_ _0210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_15_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4732_ soc.rom_encoder_0.request_data_out\[0\] _1481_ _2133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_9_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4663_ _2086_ _0172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_119_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6402_ _0275_ clknet_leaf_28_wb_clk_i soc.rom_encoder_0.request_address\[7\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3614_ _1209_ _1210_ _1211_ _1139_ _1212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_4594_ soc.spi_video_ram_1.fifo_in_address\[7\] soc.spi_video_ram_1.write_fifo.fifo_mem\[7\]\[23\]
+ _2037_ _2050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_143_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_116_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6333_ _0208_ clknet_leaf_112_wb_clk_i soc.spi_video_ram_1.buffer_index\[0\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3545_ soc.video_generator_1.v_count\[8\] soc.video_generator_1.v_count\[7\] soc.video_generator_1.v_count\[6\]
+ soc.video_generator_1.v_count\[5\] _1143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_2
XFILLER_142_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3476_ _1067_ _1066_ _1077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6264_ _0139_ clknet_leaf_98_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[7\]\[22\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_131_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5215_ _1410_ _1440_ _2473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6195_ _0075_ clknet_leaf_115_wb_clk_i soc.spi_video_ram_1.output_buffer\[5\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_97_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5146_ _2400_ _2420_ _0322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_69_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5077_ soc.spi_video_ram_1.write_fifo.fifo_mem\[3\]\[18\] soc.spi_video_ram_1.fifo_in_address\[2\]
+ _2368_ _2369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_29_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4028_ _1584_ _1585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_56_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_25_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5979_ soc.spi_video_ram_1.write_fifo.fifo_mem\[0\]\[25\] soc.spi_video_ram_1.fifo_in_address\[9\]
+ _2952_ _2980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_139_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_20_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_95_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_56_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3330_ _0875_ _0939_ _0940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_4_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5000_ _2293_ _2318_ _2319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3261_ _0853_ _0873_ _0874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_79_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3192_ _0756_ _0782_ _0793_ _0798_ _0805_ _0806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XTAP_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5902_ soc.cpu.AReg.data\[0\] _0744_ _0864_ _0930_ _2936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_5833_ net85 _2893_ _2894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_90_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_62_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5764_ _1123_ _2839_ _0847_ _2840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_50_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4715_ _2120_ _0191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5695_ soc.spi_video_ram_1.write_fifo.fifo_mem\[6\]\[1\] soc.spi_video_ram_1.fifo_in_data\[1\]
+ _2799_ _2801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4646_ soc.spi_video_ram_1.write_fifo.fifo_mem\[4\]\[18\] soc.spi_video_ram_1.fifo_in_address\[2\]
+ _2069_ _2078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_116_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4577_ _1892_ _2025_ _2041_ _0131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_143_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6316_ _0191_ clknet_leaf_145_wb_clk_i soc.spi_video_ram_1.read_value\[2\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_118_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3528_ soc.video_generator_1.v_count\[6\] _1126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_103_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3459_ _0904_ soc.cpu.ALU.x\[11\] _1061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_77_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6247_ _0122_ clknet_leaf_124_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[7\]\[5\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_130_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_57_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6178_ _0058_ clknet_leaf_114_wb_clk_i soc.spi_video_ram_1.output_buffer\[22\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_85_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5129_ _2393_ _2405_ _2406_ _2407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_57_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_67_wb_clk_i clknet_4_13_0_wb_clk_i clknet_leaf_67_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_126_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_76_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_75_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5480_ _1502_ _2594_ _2667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_8_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4500_ _1167_ _1991_ _1998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_1 net22 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4431_ _1949_ _0702_ _1950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_144_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4362_ _1710_ _1886_ _1579_ _1887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3313_ _0849_ _0923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XTAP_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6101_ _3045_ _0652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4293_ _1702_ _1818_ _1820_ _1821_ _1822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_140_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3244_ soc.cpu.AReg.data\[11\] soc.cpu.AReg.data\[10\] soc.cpu.AReg.data\[12\] soc.cpu.AReg.data\[5\]
+ _0857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XTAP_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6032_ soc.spi_video_ram_1.fifo_in_address\[4\] soc.spi_video_ram_1.write_fifo.fifo_mem\[1\]\[20\]
+ _2999_ _3009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_67_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3175_ soc.spi_video_ram_1.output_buffer\[15\] _0770_ _0789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_82_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_81_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_23_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5816_ _2318_ _2878_ _2881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_6796_ _0638_ clknet_leaf_123_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[2\]\[9\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5747_ _2827_ _0516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_136_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5678_ soc.cpu.ALU.x\[10\] _2784_ _2791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_135_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4629_ _2056_ _2069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_116_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_leaf_114_wb_clk_i clknet_4_8_0_wb_clk_i clknet_leaf_114_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_73_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_45_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_135_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput60 net60 io_out[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput71 net71 io_out[23] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_122_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput82 net82 io_out[9] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_76_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4980_ _2304_ soc.rom_encoder_0.request_address\[4\] _2287_ _2305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_51_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3931_ soc.ram_encoder_0.current_state\[2\] _1503_ _1504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_32_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3862_ _1413_ _1447_ _1448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6650_ _0492_ clknet_leaf_12_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[6\]\[2\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_20_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5601_ soc.rom_loader.writing soc.rom_loader.was_loading _2268_ _2743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_6581_ _0454_ clknet_leaf_11_wb_clk_i soc.rom_loader.rom_request vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_20_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_118_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3793_ _0779_ _0784_ _0785_ _0765_ _1379_ _1384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_5532_ soc.spi_video_ram_1.write_fifo.write_pointer\[2\] _2703_ _0698_ _2704_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_118_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5463_ soc.ram_data_out\[13\] _2604_ _2654_ _2655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_8_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5394_ soc.ram_encoder_0.initialized _1955_ _2600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_105_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4414_ _1596_ soc.spi_video_ram_1.write_fifo.fifo_mem\[6\]\[20\] _1934_ _1591_ _1935_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_114_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4345_ _1600_ soc.spi_video_ram_1.write_fifo.fifo_mem\[6\]\[13\] _1870_ _1590_ _1871_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_141_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4276_ _1756_ soc.spi_video_ram_1.write_fifo.fifo_mem\[4\]\[9\] _1805_ _1806_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6015_ _3000_ _0611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3227_ _0758_ _0836_ _0837_ _0840_ _0841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_100_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3158_ _0750_ _0771_ _0772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_27_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2019 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2008 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3089_ soc.spi_video_ram_1.start_read _0702_ _0707_ _0708_ _0709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_36_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_42_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6779_ _0621_ clknet_leaf_96_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[1\]\[21\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_7_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xcaravel_hack_soc_215 wbs_dat_o[22] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_6_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xcaravel_hack_soc_204 wbs_dat_o[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xcaravel_hack_soc_226 io_oeb[30] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_117_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1852 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1830 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1885 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1874 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1863 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_82_wb_clk_i clknet_4_9_0_wb_clk_i clknet_leaf_82_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_13_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1896 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_11_wb_clk_i clknet_4_1_0_wb_clk_i clknet_leaf_11_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_41_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4130_ soc.rom_encoder_0.output_buffer\[2\] _1671_ _1672_ soc.rom_encoder_0.request_address\[1\]
+ _1675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_69_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_68_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4061_ _1595_ soc.spi_video_ram_1.write_fifo.fifo_mem\[4\]\[18\] _1616_ _1617_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_36_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_37_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4963_ soc.rom_encoder_0.write_enable _2292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_18_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_36_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6702_ _0544_ clknet_leaf_70_wb_clk_i soc.ram_encoder_0.address\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3914_ _0676_ _1487_ _0023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4894_ soc.rom_encoder_0.input_buffer\[3\] _2249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6633_ _0475_ net89 soc.cpu.ALU.x\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_60_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3845_ _1410_ _1431_ _1432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_20_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6564_ _0437_ clknet_leaf_73_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[5\]\[12\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3776_ _0808_ _0822_ _1364_ _1367_ _1368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_6495_ _0368_ clknet_leaf_43_wb_clk_i soc.ram_encoder_0.request_data_out\[8\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5515_ soc.hack_clock_0.counter\[0\] soc.hack_clock_0.counter\[1\] _2693_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__and2_1
X_5446_ _2516_ _2624_ _2625_ _2641_ _2642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_5377_ _2587_ _0386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_59_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4328_ _1854_ _0069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4259_ soc.spi_video_ram_1.write_fifo.fifo_mem\[7\]\[8\] _1790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_101_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_124_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_77_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_66_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_74_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1693 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3630_ _1225_ _1227_ _1228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_3561_ soc.boot_loading_offset\[1\] _1144_ _1159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_128_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5300_ _2537_ _2538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_3492_ _0845_ _0887_ soc.cpu.AReg.data\[12\] _0880_ _1093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_6280_ _0155_ clknet_leaf_82_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[4\]\[9\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_6_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5231_ soc.rom_encoder_0.initializing_step\[4\] _2484_ _2485_ _2486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_45_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5162_ _2400_ _2432_ _0326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_64_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4113_ _1120_ _1660_ _1661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_69_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5093_ soc.spi_video_ram_1.write_fifo.fifo_mem\[3\]\[26\] soc.spi_video_ram_1.fifo_in_address\[10\]
+ _2368_ _2377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_112_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4044_ _1600_ _1601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_80_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5995_ soc.spi_video_ram_1.fifo_in_data\[2\] soc.spi_video_ram_1.write_fifo.fifo_mem\[1\]\[2\]
+ _2986_ _2990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_24_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4946_ soc.rom_encoder_0.data_out\[8\] soc.rom_encoder_0.request_data_out\[8\] _2276_
+ _2283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4877_ _2226_ _2234_ _2237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6616_ _0473_ clknet_leaf_72_wb_clk_i net83 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3828_ soc.rom_encoder_0.output_bits_left\[3\] _1415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_21_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6547_ _0420_ clknet_leaf_31_wb_clk_i soc.hack_clock_0.counter\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_116_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3759_ _1189_ _1195_ _1351_ _1356_ _1357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_118_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6478_ _0351_ clknet_leaf_45_wb_clk_i soc.ram_encoder_0.input_buffer\[4\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_134_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5429_ soc.ram_encoder_0.request_data_out\[5\] _2606_ _2629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_48_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_120_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_4_0_0_wb_clk_i clknet_0_wb_clk_i clknet_4_0_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_34_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2180 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4800_ _0759_ _2186_ _2187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5780_ soc.cpu.PC.REG.data\[2\] _2853_ _2854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_34_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4731_ _1671_ _2130_ _2131_ _2132_ _0195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4662_ soc.spi_video_ram_1.write_fifo.fifo_mem\[4\]\[26\] soc.spi_video_ram_1.fifo_in_address\[10\]
+ _2057_ _2086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6401_ _0274_ clknet_leaf_28_wb_clk_i soc.rom_encoder_0.request_address\[6\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3613_ _1142_ _1143_ _1211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_134_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4593_ _2049_ _0139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6332_ _0207_ clknet_leaf_24_wb_clk_i soc.rom_encoder_0.output_buffer\[19\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3544_ soc.video_generator_1.v_count\[9\] _1142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_135_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_116_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3475_ _1072_ _1075_ _1076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6263_ _0138_ clknet_leaf_95_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[7\]\[21\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_143_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5214_ soc.rom_encoder_0.initializing_step\[1\] _1438_ _2472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6194_ _0074_ clknet_leaf_113_wb_clk_i soc.spi_video_ram_1.output_buffer\[6\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_111_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5145_ soc.cpu.instruction\[5\] _2392_ _2419_ _2420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_84_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5076_ _2216_ _2368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_4027_ _1583_ _1584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_25_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5978_ _2979_ _0595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4929_ soc.rom_encoder_0.data_out\[0\] soc.rom_encoder_0.request_data_out\[0\] _2272_
+ _2274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xclkbuf_leaf_139_wb_clk_i clknet_4_2_0_wb_clk_i clknet_leaf_139_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_60_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_112_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3260_ _0854_ _0855_ _0863_ _0872_ soc.cpu.ALU.zy _0873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_79_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3191_ soc.spi_video_ram_1.buffer_index\[4\] _0780_ _0804_ _0805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_120_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5901_ _2934_ _2932_ _2935_ _0562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_19_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_35_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5832_ _2688_ _2689_ _2692_ _2893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_62_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5763_ _1069_ _1108_ _2838_ _2839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_4714_ net11 soc.spi_video_ram_1.read_value\[2\] _2117_ _2120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5694_ _2800_ _0490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_30_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4645_ _2077_ _0163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4576_ soc.spi_video_ram_1.fifo_in_data\[14\] _2026_ _2041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_115_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6315_ _0190_ clknet_leaf_144_wb_clk_i soc.spi_video_ram_1.read_value\[1\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3527_ soc.video_generator_1.v_count\[9\] _1125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_3
XFILLER_143_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_131_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3458_ _1042_ _1045_ _1055_ _0972_ _1060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_6246_ _0121_ clknet_leaf_125_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[7\]\[4\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_97_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3389_ soc.ram_data_out\[7\] _0869_ _0868_ net44 _0854_ _0995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_85_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6177_ _0057_ clknet_leaf_134_wb_clk_i soc.spi_video_ram_1.output_buffer\[23\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5128_ net7 _2223_ _2406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5059_ _2359_ _0296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_111_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_107_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_36_wb_clk_i clknet_4_7_0_wb_clk_i clknet_leaf_36_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_121_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_32_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_2 net25 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4430_ soc.spi_video_ram_1.fifo_read_request _1949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_144_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_99_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6100_ soc.spi_video_ram_1.write_fifo.fifo_mem\[2\]\[23\] soc.spi_video_ram_1.fifo_in_address\[7\]
+ _3019_ _3045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4361_ soc.spi_video_ram_1.write_fifo.fifo_mem\[2\]\[14\] soc.spi_video_ram_1.write_fifo.fifo_mem\[3\]\[14\]
+ _1582_ _1886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_101_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3312_ soc.cpu.ALU.no _0922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XTAP_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4292_ _0703_ _1608_ _1821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_100_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3243_ soc.cpu.AReg.data\[4\] soc.cpu.AReg.data\[7\] soc.cpu.AReg.data\[6\] _0856_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_79_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6031_ _3008_ _0619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3174_ _0783_ soc.spi_video_ram_1.output_buffer\[14\] _0788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_39_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_63_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5815_ _2847_ _2879_ _2880_ _2849_ _0530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_22_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6795_ _0637_ clknet_leaf_115_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[2\]\[8\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_22_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5746_ soc.spi_video_ram_1.write_fifo.fifo_mem\[6\]\[26\] soc.spi_video_ram_1.fifo_in_address\[10\]
+ _2798_ _2827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5677_ _1039_ _2778_ _2790_ _0483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4628_ _2068_ _0155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_123_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4559_ soc.spi_video_ram_1.fifo_in_data\[6\] _2026_ _2032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_104_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_103_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6229_ _0104_ clknet_leaf_15_wb_clk_i soc.spi_video_ram_1.fifo_in_data\[3\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_58_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput61 net61 io_out[13] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput50 net50 io_oeb[16] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput72 net72 io_out[24] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_122_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput83 net83 la_data_out[27] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_68_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3930_ soc.ram_encoder_0.current_state\[1\] _1502_ _1503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_63_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3861_ soc.rom_encoder_0.output_buffer\[18\] _1417_ _1442_ soc.rom_encoder_0.request_data_out\[14\]
+ _1447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_32_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5600_ soc.rom_loader.rom_request _2458_ soc.rom_loader.writing _2742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3792_ soc.spi_video_ram_1.buffer_index\[4\] _1382_ _1383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_6580_ _0453_ clknet_leaf_109_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[5\]\[28\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_75_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5531_ _0694_ _2703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_118_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5462_ _2524_ _2624_ _2625_ _2653_ _2654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_5393_ soc.ram_encoder_0.initializing_step\[0\] _2596_ _2598_ _2599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_99_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4413_ _1756_ _1933_ _1934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4344_ _1755_ _1869_ _1870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_140_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_143_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4275_ _1593_ _1804_ _1586_ _1805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_6014_ soc.spi_video_ram_1.fifo_in_data\[11\] soc.spi_video_ram_1.write_fifo.fifo_mem\[1\]\[11\]
+ _2999_ _3000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_86_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3226_ _0760_ _0838_ _0839_ _0811_ soc.spi_video_ram_1.buffer_index\[4\] _0840_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_82_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3157_ soc.spi_video_ram_1.buffer_index\[1\] _0770_ _0771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_39_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2009 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3088_ soc.spi_video_ram_1.current_state\[2\] _0708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_36_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_42_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xclkbuf_4_13_0_wb_clk_i clknet_0_wb_clk_i clknet_4_13_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_51_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_11_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6778_ _0620_ clknet_leaf_88_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[1\]\[20\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5729_ _2818_ _0507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_10_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xcaravel_hack_soc_205 wbs_dat_o[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_136_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xcaravel_hack_soc_227 io_oeb[31] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
Xcaravel_hack_soc_216 wbs_dat_o[23] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_132_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_73_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_100_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1842 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1820 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1831 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1875 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1864 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1853 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1897 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1886 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_51_wb_clk_i clknet_4_6_0_wb_clk_i clknet_leaf_51_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_54_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_6_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4060_ _1596_ _1615_ _1616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_110_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4962_ _2291_ _0267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_51_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6701_ _0543_ clknet_leaf_70_wb_clk_i soc.ram_encoder_0.address\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4893_ _2247_ _2242_ _2248_ _0241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_33_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3913_ _1430_ _1485_ _1486_ net64 _1487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_6632_ _0474_ net89 soc.cpu.ALU.x\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3844_ _1430_ _1431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_20_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_20_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6563_ _0436_ clknet_leaf_94_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[5\]\[11\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_9_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3775_ _1365_ _1366_ _1367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_118_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6494_ _0367_ clknet_leaf_61_wb_clk_i soc.ram_encoder_0.request_data_out\[7\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5514_ soc.hack_clock_0.counter\[0\] soc.hack_clock_0.counter\[1\] _2692_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5445_ soc.ram_encoder_0.request_data_out\[9\] _2605_ _2641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_114_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5376_ soc.ram_encoder_0.address\[10\] soc.ram_encoder_0.request_address\[10\] _2581_
+ _2587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_141_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4327_ soc.spi_video_ram_1.output_buffer\[11\] _1612_ _1825_ _1853_ _1854_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_102_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4258_ _1585_ _1787_ _1788_ _1710_ _1789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_74_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3209_ _0760_ _0822_ _0823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_41_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4189_ soc.spi_video_ram_1.write_fifo.fifo_mem\[4\]\[3\] soc.spi_video_ram_1.write_fifo.fifo_mem\[5\]\[3\]
+ soc.spi_video_ram_1.write_fifo.fifo_mem\[6\]\[3\] soc.spi_video_ram_1.write_fifo.fifo_mem\[7\]\[3\]
+ _1724_ _1587_ _1725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_27_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_11_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xcaravel_hack_soc_92 io_oeb[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_73_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_33_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1694 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_42_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3560_ soc.boot_loading_offset\[0\] _1140_ _1158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_3491_ _0990_ _1091_ _1092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_5230_ _2221_ _2380_ _2485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_64_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5161_ _1011_ _2392_ _2431_ _2432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_68_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_84_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4112_ _0954_ _1659_ _1660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5092_ _2376_ _0312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_56_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4043_ _1583_ _1600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_83_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5994_ _1698_ _2988_ _2989_ _0601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4945_ _2282_ _0259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_80_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4876_ _2222_ _2231_ _2236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_20_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3827_ soc.rom_encoder_0.output_bits_left\[4\] _1414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6615_ _0472_ clknet_leaf_6_wb_clk_i soc.rom_loader.wait_fall_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_119_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6546_ _0419_ clknet_leaf_31_wb_clk_i soc.hack_clock_0.counter\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3758_ _1352_ _1355_ _1356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_6477_ _0350_ clknet_leaf_45_wb_clk_i soc.ram_encoder_0.input_buffer\[3\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3689_ _1196_ _1281_ _1287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_121_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5428_ _2615_ _2628_ _0396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_121_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5359_ soc.ram_encoder_0.address\[2\] soc.ram_encoder_0.request_address\[2\] _2566_
+ _2578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_58_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_70_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2170 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2181 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4730_ soc.rom_encoder_0.request_address\[6\] _1672_ _2132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4661_ _2085_ _0171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6400_ _0273_ clknet_leaf_32_wb_clk_i soc.rom_encoder_0.request_address\[5\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3612_ _1163_ _1165_ _1169_ _1170_ _1210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_128_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6331_ _0206_ clknet_leaf_24_wb_clk_i soc.rom_encoder_0.output_buffer\[18\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_31_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4592_ soc.spi_video_ram_1.fifo_in_address\[6\] soc.spi_video_ram_1.write_fifo.fifo_mem\[7\]\[22\]
+ _2037_ _2049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_3543_ soc.boot_loading_offset\[0\] _1140_ _1141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_143_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_3474_ _0926_ _1074_ _1075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_6_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6262_ _0137_ clknet_leaf_119_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[7\]\[20\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_142_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5213_ _1438_ _2380_ _2382_ _2471_ _0338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_6193_ _0073_ clknet_leaf_114_wb_clk_i soc.spi_video_ram_1.output_buffer\[7\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5144_ _2245_ _2413_ _2414_ _2418_ _2419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_9_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5075_ _2367_ _0304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_57_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4026_ _1582_ _1583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_65_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5977_ soc.spi_video_ram_1.write_fifo.fifo_mem\[0\]\[24\] soc.spi_video_ram_1.fifo_in_address\[8\]
+ _2952_ _2979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4928_ _2089_ _2272_ _2273_ _0251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_121_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4859_ _2220_ _0235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_5_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6529_ _0402_ clknet_leaf_57_wb_clk_i soc.ram_data_out\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_leaf_108_wb_clk_i clknet_4_10_0_wb_clk_i clknet_leaf_108_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_134_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_12_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_137_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3190_ _0762_ _0803_ _0804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_39_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5900_ _0741_ _2935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_34_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5831_ _2847_ _2891_ _2892_ _0743_ _0534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_5762_ _2832_ _2833_ _2834_ _2837_ _2838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_22_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_6_wb_clk_i clknet_4_1_0_wb_clk_i clknet_leaf_6_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_4713_ _1349_ _2117_ _2119_ _0190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5693_ soc.spi_video_ram_1.write_fifo.fifo_mem\[6\]\[0\] soc.spi_video_ram_1.fifo_in_data\[0\]
+ _2799_ _2800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4644_ soc.spi_video_ram_1.write_fifo.fifo_mem\[4\]\[17\] soc.spi_video_ram_1.fifo_in_address\[1\]
+ _2069_ _2077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_129_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4575_ _1869_ _2025_ _2040_ _0130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_144_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3526_ _0883_ _1123_ _1124_ soc.cpu.PC.in\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_6314_ _0189_ clknet_leaf_144_wb_clk_i soc.spi_video_ram_1.read_value\[0\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_143_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6245_ _0120_ clknet_leaf_14_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[7\]\[3\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_143_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3457_ _0883_ _1058_ _1059_ soc.cpu.PC.in\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_6176_ _0056_ clknet_leaf_64_wb_clk_i soc.ram_encoder_0.output_buffer\[1\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3388_ _0849_ _0993_ _0994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_5127_ soc.rom_encoder_0.request_data_out\[2\] _2395_ _2405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_58_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_84_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5058_ soc.spi_video_ram_1.write_fifo.fifo_mem\[3\]\[9\] soc.spi_video_ram_1.fifo_in_data\[9\]
+ _2357_ _2359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_29_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4009_ soc.ram_encoder_0.output_buffer\[14\] _1555_ _1530_ soc.ram_encoder_0.request_data_out\[10\]
+ _1559_ _1569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_85_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_122_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_76_wb_clk_i clknet_4_15_0_wb_clk_i clknet_leaf_76_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_76_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_21_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_3 net72 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4360_ _1756_ soc.spi_video_ram_1.write_fifo.fifo_mem\[0\]\[14\] _1884_ _1885_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_141_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3311_ _0884_ _0920_ _0921_ soc.cpu.PC.in\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_112_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4291_ _1580_ _1819_ _1820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_113_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3242_ soc.cpu.AReg.data\[0\] _0855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_2
X_6030_ soc.spi_video_ram_1.fifo_in_address\[3\] soc.spi_video_ram_1.write_fifo.fifo_mem\[1\]\[19\]
+ _2999_ _3008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3173_ _0776_ soc.spi_video_ram_1.output_buffer\[12\] _0772_ soc.spi_video_ram_1.output_buffer\[13\]
+ _0787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_20_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_39_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_67_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_35_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_63_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5814_ soc.cpu.PC.in\[10\] _2851_ _2880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_23_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6794_ _0636_ clknet_leaf_127_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[2\]\[7\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5745_ _2826_ _0515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_22_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5676_ soc.cpu.ALU.x\[9\] _2784_ _2790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_135_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4627_ soc.spi_video_ram_1.write_fifo.fifo_mem\[4\]\[9\] soc.spi_video_ram_1.fifo_in_data\[9\]
+ _2058_ _2068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_117_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_116_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4558_ _1743_ _2025_ _2031_ _0122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_143_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3509_ _0845_ soc.cpu.instruction\[13\] soc.cpu.AReg.data\[13\] _0880_ _1109_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_4489_ soc.video_generator_1.v_count\[3\] _1989_ _1991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_89_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6228_ _0103_ clknet_leaf_16_wb_clk_i soc.spi_video_ram_1.fifo_in_data\[2\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_44_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_131_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6159_ _0039_ clknet_leaf_117_wb_clk_i soc.spi_video_ram_1.output_buffer\[1\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_66_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_26_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xclkbuf_leaf_123_wb_clk_i clknet_4_9_0_wb_clk_i clknet_leaf_123_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_40_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_108_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput51 net51 io_oeb[17] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_110_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput62 net62 io_out[14] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput73 net73 io_out[25] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_110_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3860_ _1432_ _1445_ _1446_ _0676_ _0010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_3791_ _0763_ _0753_ _1382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_31_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5530_ _2691_ _2702_ _0424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XPHY_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5461_ soc.ram_encoder_0.request_data_out\[13\] _2605_ _2653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_68_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4412_ soc.spi_video_ram_1.write_fifo.fifo_mem\[7\]\[20\] _1933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5392_ soc.ram_encoder_0.initializing_step\[0\] _2597_ _2598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_113_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4343_ soc.spi_video_ram_1.write_fifo.fifo_mem\[7\]\[13\] _1869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4274_ soc.spi_video_ram_1.write_fifo.fifo_mem\[5\]\[9\] _1804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_101_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3225_ soc.spi_video_ram_1.output_buffer\[2\] soc.spi_video_ram_1.output_buffer\[3\]
+ _0750_ _0839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6013_ _2985_ _2999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_86_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3156_ _0749_ _0769_ _0753_ _0770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_54_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3087_ _0702_ _0706_ soc.spi_video_ram_1.initialized _0707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_82_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6777_ _0619_ clknet_leaf_89_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[1\]\[19\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_22_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3989_ soc.ram_encoder_0.output_buffer\[11\] _1519_ _1552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_109_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5728_ soc.spi_video_ram_1.write_fifo.fifo_mem\[6\]\[17\] soc.spi_video_ram_1.fifo_in_address\[1\]
+ _2810_ _2818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xcaravel_hack_soc_206 wbs_dat_o[13] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_109_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5659_ soc.cpu.ALU.x\[1\] _2779_ _2781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xcaravel_hack_soc_217 wbs_dat_o[24] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xcaravel_hack_soc_228 io_oeb[32] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_105_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_78_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_77_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1843 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1821 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1832 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1810 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1865 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1854 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_42_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1898 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1887 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_142_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_91_wb_clk_i clknet_4_14_0_wb_clk_i clknet_leaf_91_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_111_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xclkbuf_leaf_20_wb_clk_i clknet_4_4_0_wb_clk_i clknet_leaf_20_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_1_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_36_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4961_ soc.rom_encoder_0.data_out\[15\] soc.rom_encoder_0.request_data_out\[15\]
+ _2287_ _2291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_45_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6700_ _0542_ clknet_leaf_70_wb_clk_i soc.ram_encoder_0.address\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4892_ net7 _2243_ _1955_ _2248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3912_ soc.rom_encoder_0.initializing_step\[4\] soc.rom_encoder_0.initializing_step\[3\]
+ _1430_ _1432_ _1486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_6631_ soc.cpu.PC.in\[14\] net88 soc.cpu.AReg.data\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_60_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3843_ _1424_ _1429_ _1430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_32_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6562_ _0435_ clknet_leaf_90_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[5\]\[10\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3774_ _0811_ _0825_ _0827_ _0815_ _1366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_121_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6493_ _0366_ clknet_leaf_63_wb_clk_i soc.ram_encoder_0.request_data_out\[6\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5513_ soc.hack_clock_0.counter\[0\] _2691_ _0418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5444_ _2615_ _2640_ _0400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5375_ _2586_ _0385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_114_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_101_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4326_ _1821_ _1844_ _1849_ _1850_ _1852_ _1853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_101_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4257_ _1600_ soc.spi_video_ram_1.write_fifo.fifo_mem\[4\]\[8\] _1788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_86_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4188_ _1583_ _1724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_3208_ _0776_ _0820_ _0821_ _0822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3139_ soc.spi_video_ram_1.buffer_index\[2\] _0752_ _0753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_28_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_51_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6829_ _0671_ clknet_leaf_50_wb_clk_i soc.ram_encoder_0.data_out\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_51_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_74_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xcaravel_hack_soc_93 io_oeb[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_18_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_105_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1695 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3490_ _0954_ _1076_ _1087_ _1090_ _1091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XFILLER_10_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5160_ _2254_ _2413_ _2414_ _2430_ _2431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_4111_ _1111_ _1114_ _1659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5091_ soc.spi_video_ram_1.write_fifo.fifo_mem\[3\]\[25\] soc.spi_video_ram_1.fifo_in_address\[9\]
+ _2368_ _2376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_110_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4042_ _1595_ soc.spi_video_ram_1.write_fifo.fifo_mem\[4\]\[16\] _1598_ _1599_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_49_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5993_ soc.spi_video_ram_1.fifo_in_data\[1\] _2988_ _2989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4944_ soc.rom_encoder_0.data_out\[7\] soc.rom_encoder_0.request_data_out\[7\] _2276_
+ _2282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_80_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4875_ _2233_ _2235_ _0236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6614_ _0471_ clknet_leaf_20_wb_clk_i soc.rom_loader.current_address\[14\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3826_ _1406_ _1412_ _1413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_118_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6545_ _0418_ clknet_leaf_31_wb_clk_i soc.hack_clock_0.counter\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3757_ _1353_ _1354_ _1355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_118_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6476_ _0349_ clknet_leaf_58_wb_clk_i soc.ram_encoder_0.input_buffer\[2\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3688_ _1215_ _1220_ _1286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_133_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5427_ soc.ram_data_out\[4\] _2603_ _2627_ _2628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_114_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5358_ _2577_ _0377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_87_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4309_ _0729_ _1354_ _1836_ _1837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_5289_ soc.ram_encoder_0.input_buffer\[11\] _2528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_102_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_79_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_80_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2171 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2160 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2182 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4660_ soc.spi_video_ram_1.write_fifo.fifo_mem\[4\]\[25\] soc.spi_video_ram_1.fifo_in_address\[9\]
+ _2057_ _2085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_30_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3611_ soc.boot_loading_offset\[0\] _1209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6330_ _0205_ clknet_leaf_24_wb_clk_i soc.rom_encoder_0.output_buffer\[17\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4591_ _2048_ _0138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_50_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3542_ _1125_ _1139_ _1128_ _1140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_115_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3473_ _1011_ _1073_ _1074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6261_ _0136_ clknet_leaf_118_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[7\]\[19\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_97_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6192_ _0072_ clknet_leaf_110_wb_clk_i soc.spi_video_ram_1.output_buffer\[8\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_5212_ _0689_ _2471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_5143_ soc.rom_encoder_0.request_data_out\[5\] _2395_ _2418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5074_ soc.spi_video_ram_1.write_fifo.fifo_mem\[3\]\[17\] soc.spi_video_ram_1.fifo_in_address\[1\]
+ _2357_ _2367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_56_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4025_ _0000_ _1582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_53_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5976_ _2978_ _0594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4927_ soc.rom_encoder_0.request_write _2272_ _2273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_60_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4858_ _1955_ _1956_ _2220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_3809_ soc.spi_video_ram_1.buffer_index\[4\] _1382_ soc.spi_video_ram_1.buffer_index\[5\]
+ _1400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_20_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4789_ _0776_ _2177_ _2178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_20_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6528_ _0401_ clknet_leaf_57_wb_clk_i soc.ram_data_out\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_107_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6459_ _0332_ clknet_leaf_19_wb_clk_i soc.cpu.instruction\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_134_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_75_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_29_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5830_ soc.cpu.PC.in\[14\] _2851_ _2892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_61_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5761_ _0989_ _1024_ _2836_ _2837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_50_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4712_ net10 _2117_ _2119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5692_ _2798_ _2799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_4643_ _2076_ _0162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_30_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4574_ soc.spi_video_ram_1.fifo_in_data\[13\] _2026_ _2040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_104_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3525_ _0845_ soc.cpu.instruction\[14\] soc.cpu.AReg.data\[14\] _0880_ _1124_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_6313_ _0188_ clknet_leaf_141_wb_clk_i net68 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6244_ _0119_ clknet_leaf_12_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[7\]\[2\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_3456_ _0845_ _0923_ soc.cpu.AReg.data\[10\] _0880_ _1059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_6175_ _0055_ clknet_leaf_66_wb_clk_i soc.ram_encoder_0.output_buffer\[2\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_85_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3387_ _0904_ soc.cpu.ALU.x\[7\] _0993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_130_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5126_ _2400_ _2404_ _0318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_57_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5057_ _2358_ _0295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_38_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4008_ _1522_ _1567_ _1568_ _0036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_26_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_26_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5959_ soc.spi_video_ram_1.write_fifo.fifo_mem\[0\]\[15\] soc.spi_video_ram_1.fifo_in_data\[15\]
+ _2964_ _2970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_40_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_leaf_45_wb_clk_i clknet_4_7_0_wb_clk_i clknet_leaf_45_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_43_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_4 net81 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3310_ _0846_ soc.cpu.DMuxJMP.sel\[2\] soc.cpu.AReg.data\[2\] _0881_ _0921_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_125_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4290_ soc.spi_video_ram_1.write_fifo.fifo_mem\[0\]\[10\] soc.spi_video_ram_1.write_fifo.fifo_mem\[1\]\[10\]
+ soc.spi_video_ram_1.write_fifo.fifo_mem\[2\]\[10\] soc.spi_video_ram_1.write_fifo.fifo_mem\[3\]\[10\]
+ _1583_ _1586_ _1819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_141_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3241_ soc.cpu.instruction\[12\] _0854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_67_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3172_ _0784_ _0785_ _0775_ _0786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_26_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5813_ soc.cpu.PC.REG.data\[10\] _2878_ _2879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_6793_ _0635_ clknet_leaf_123_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[2\]\[6\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_50_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5744_ soc.spi_video_ram_1.write_fifo.fifo_mem\[6\]\[25\] soc.spi_video_ram_1.fifo_in_address\[9\]
+ _2798_ _2826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5675_ _1024_ _2778_ _2789_ _0482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_129_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4626_ _2067_ _0154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_144_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4557_ soc.spi_video_ram_1.fifo_in_data\[5\] _2026_ _2031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_104_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3508_ _0990_ _1107_ _1108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_4488_ soc.video_generator_1.v_count\[3\] _1989_ _1990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_106_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3439_ _0923_ _1041_ _1042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_6227_ _0102_ clknet_leaf_52_wb_clk_i soc.spi_video_ram_1.fifo_in_data\[1\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_131_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6158_ _0038_ clknet_leaf_60_wb_clk_i soc.ram_encoder_0.output_buffer\[19\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_98_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5109_ _2223_ _2228_ _2388_ _2389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_46_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6089_ _3039_ _0646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_85_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_26_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_25_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xoutput52 net52 io_oeb[18] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_107_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput63 net63 io_out[15] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_123_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput74 net74 io_out[27] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_110_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3790_ _0775_ _0787_ _1379_ _1380_ _1381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_20_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_5460_ _2471_ _2652_ _0404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_133_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4411_ _1601_ soc.spi_video_ram_1.write_fifo.fifo_mem\[4\]\[20\] _1931_ _1932_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5391_ _1405_ _2334_ _2597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4342_ _1756_ soc.spi_video_ram_1.write_fifo.fifo_mem\[4\]\[13\] _1867_ _1868_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4273_ soc.spi_video_ram_1.write_fifo.fifo_mem\[6\]\[9\] soc.spi_video_ram_1.write_fifo.fifo_mem\[7\]\[9\]
+ _1584_ _1803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_28_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6012_ _2998_ _0610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3224_ soc.spi_video_ram_1.output_buffer\[6\] soc.spi_video_ram_1.output_buffer\[7\]
+ _0750_ _0838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
.ends

