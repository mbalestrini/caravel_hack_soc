VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO caravel_hack_soc
  CLASS BLOCK ;
  FOREIGN caravel_hack_soc ;
  ORIGIN 0.000 0.000 ;
  SIZE 1000.000 BY 1000.000 ;
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 346.080 4.000 346.640 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 460.320 4.000 460.880 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 413.280 4.000 413.840 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 964.320 996.000 964.880 999.000 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 356.160 4.000 356.720 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 551.040 996.000 551.600 999.000 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 194.880 999.000 195.440 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 288.960 1.000 289.520 4.000 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 221.760 996.000 222.320 999.000 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 443.520 4.000 444.080 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 994.560 999.000 995.120 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 803.040 996.000 803.600 999.000 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 581.280 996.000 581.840 999.000 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 947.520 996.000 948.080 999.000 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 20.160 996.000 20.720 999.000 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 134.400 1.000 134.960 4.000 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 127.680 996.000 128.240 999.000 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 164.640 996.000 165.200 999.000 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 107.520 999.000 108.080 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 238.560 4.000 239.120 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 40.320 996.000 40.880 999.000 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 974.400 999.000 974.960 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 104.160 4.000 104.720 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 702.240 1.000 702.800 4.000 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 144.480 996.000 145.040 999.000 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 598.080 1.000 598.640 4.000 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 981.120 4.000 981.680 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 897.120 996.000 897.680 999.000 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 211.680 996.000 212.240 999.000 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 258.720 4.000 259.280 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 164.640 999.000 165.200 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 423.360 4.000 423.920 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 897.120 1.000 897.680 4.000 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 974.400 4.000 974.960 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 228.480 4.000 229.040 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 262.080 999.000 262.640 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 974.400 1.000 974.960 4.000 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 850.080 996.000 850.640 999.000 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 30.240 996.000 30.800 999.000 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 682.080 4.000 682.640 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 624.960 4.000 625.520 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 752.640 4.000 753.200 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 856.800 1.000 857.360 4.000 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 981.120 1.000 981.680 4.000 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 530.880 996.000 531.440 999.000 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 577.920 4.000 578.480 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 97.440 996.000 98.000 999.000 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 789.600 4.000 790.160 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 403.200 1.000 403.760 4.000 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 77.280 999.000 77.840 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 846.720 1.000 847.280 4.000 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 94.080 1.000 94.640 4.000 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 252.000 999.000 252.560 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 94.080 4.000 94.640 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 221.760 999.000 222.320 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 356.160 1.000 356.720 4.000 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 829.920 1.000 830.480 4.000 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 665.280 4.000 665.840 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 934.080 4.000 934.640 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 204.960 996.000 205.520 999.000 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 645.120 1.000 645.680 4.000 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 36.960 4.000 37.520 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 695.520 999.000 696.080 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 154.560 999.000 155.120 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 819.840 4.000 820.400 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 383.040 4.000 383.600 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 561.120 996.000 561.680 999.000 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 934.080 1.000 934.640 4.000 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 836.640 4.000 837.200 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 339.360 999.000 339.920 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 996.000 0.560 999.000 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 964.320 999.000 964.880 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 483.840 996.000 484.400 999.000 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 57.120 999.000 57.680 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 406.560 999.000 407.120 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 396.480 999.000 397.040 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 191.520 4.000 192.080 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 974.400 996.000 974.960 999.000 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 880.320 999.000 880.880 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 984.480 999.000 985.040 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 742.560 4.000 743.120 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 393.120 1.000 393.680 4.000 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 829.920 999.000 830.480 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 114.240 1.000 114.800 4.000 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 836.640 1.000 837.200 4.000 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 655.200 1.000 655.760 4.000 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 67.200 1.000 67.760 4.000 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 682.080 1.000 682.640 4.000 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 450.240 1.000 450.800 4.000 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 336.000 1.000 336.560 4.000 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 134.400 4.000 134.960 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 735.840 996.000 736.400 999.000 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 463.680 996.000 464.240 999.000 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 423.360 1.000 423.920 4.000 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 705.600 996.000 706.160 999.000 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 742.560 1.000 743.120 4.000 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 638.400 996.000 638.960 999.000 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 944.160 1.000 944.720 4.000 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 917.280 996.000 917.840 999.000 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 211.680 999.000 212.240 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 840.000 996.000 840.560 999.000 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 319.200 999.000 319.760 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 665.280 1.000 665.840 4.000 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 648.480 999.000 649.040 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 238.560 1.000 239.120 4.000 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 937.440 999.000 938.000 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 927.360 999.000 927.920 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 715.680 999.000 716.240 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 26.880 4.000 27.440 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 47.040 4.000 47.600 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 567.840 4.000 568.400 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 628.320 996.000 628.880 999.000 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 258.720 1.000 259.280 4.000 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 510.720 4.000 511.280 ;
    END
  END io_out[9]
  PIN irq[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 702.240 4.000 702.800 ;
    END
  END irq[0]
  PIN irq[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 403.200 4.000 403.760 ;
    END
  END irq[1]
  PIN irq[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 305.760 1.000 306.320 4.000 ;
    END
  END irq[2]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 406.560 996.000 407.120 999.000 ;
    END
  END la_data_in[0]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 937.440 996.000 938.000 999.000 ;
    END
  END la_data_in[10]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 470.400 1.000 470.960 4.000 ;
    END
  END la_data_in[11]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 604.800 4.000 605.360 ;
    END
  END la_data_in[12]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 144.480 999.000 145.040 ;
    END
  END la_data_in[13]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 366.240 999.000 366.800 ;
    END
  END la_data_in[14]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 692.160 4.000 692.720 ;
    END
  END la_data_in[15]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 231.840 996.000 232.400 999.000 ;
    END
  END la_data_in[16]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 204.960 999.000 205.520 ;
    END
  END la_data_in[17]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 752.640 999.000 753.200 ;
    END
  END la_data_in[18]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 443.520 999.000 444.080 ;
    END
  END la_data_in[19]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 762.720 996.000 763.280 999.000 ;
    END
  END la_data_in[1]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 510.720 996.000 511.280 999.000 ;
    END
  END la_data_in[20]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 161.280 4.000 161.840 ;
    END
  END la_data_in[21]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 618.240 996.000 618.800 999.000 ;
    END
  END la_data_in[22]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 903.840 4.000 904.400 ;
    END
  END la_data_in[23]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 433.440 996.000 434.000 999.000 ;
    END
  END la_data_in[24]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 241.920 999.000 242.480 ;
    END
  END la_data_in[25]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 325.920 1.000 326.480 4.000 ;
    END
  END la_data_in[26]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 73.920 4.000 74.480 ;
    END
  END la_data_in[27]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 366.240 4.000 366.800 ;
    END
  END la_data_in[28]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 759.360 4.000 759.920 ;
    END
  END la_data_in[29]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 675.360 4.000 675.920 ;
    END
  END la_data_in[2]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 77.280 996.000 77.840 999.000 ;
    END
  END la_data_in[30]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 887.040 4.000 887.600 ;
    END
  END la_data_in[31]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 504.000 996.000 504.560 999.000 ;
    END
  END la_data_in[32]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 850.080 999.000 850.640 ;
    END
  END la_data_in[33]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 309.120 996.000 309.680 999.000 ;
    END
  END la_data_in[34]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 416.640 996.000 417.200 999.000 ;
    END
  END la_data_in[35]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 540.960 999.000 541.520 ;
    END
  END la_data_in[36]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 346.080 1.000 346.640 4.000 ;
    END
  END la_data_in[37]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 480.480 1.000 481.040 4.000 ;
    END
  END la_data_in[38]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 336.000 4.000 336.560 ;
    END
  END la_data_in[39]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 618.240 999.000 618.800 ;
    END
  END la_data_in[3]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 10.080 999.000 10.640 ;
    END
  END la_data_in[40]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 944.160 4.000 944.720 ;
    END
  END la_data_in[41]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 725.760 999.000 726.320 ;
    END
  END la_data_in[42]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 614.880 1.000 615.440 4.000 ;
    END
  END la_data_in[43]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 473.760 996.000 474.320 999.000 ;
    END
  END la_data_in[44]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 134.400 996.000 134.960 999.000 ;
    END
  END la_data_in[45]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 87.360 996.000 87.920 999.000 ;
    END
  END la_data_in[46]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 396.480 996.000 397.040 999.000 ;
    END
  END la_data_in[47]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 460.320 1.000 460.880 4.000 ;
    END
  END la_data_in[48]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 520.800 4.000 521.360 ;
    END
  END la_data_in[49]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 819.840 996.000 820.400 999.000 ;
    END
  END la_data_in[4]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 305.760 4.000 306.320 ;
    END
  END la_data_in[50]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 268.800 4.000 269.360 ;
    END
  END la_data_in[51]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 299.040 4.000 299.600 ;
    END
  END la_data_in[52]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 30.240 999.000 30.800 ;
    END
  END la_data_in[53]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 366.240 1.000 366.800 4.000 ;
    END
  END la_data_in[54]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 907.200 999.000 907.760 ;
    END
  END la_data_in[55]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 171.360 1.000 171.920 4.000 ;
    END
  END la_data_in[56]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 262.080 996.000 262.640 999.000 ;
    END
  END la_data_in[57]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 376.320 996.000 376.880 999.000 ;
    END
  END la_data_in[58]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 588.000 1.000 588.560 4.000 ;
    END
  END la_data_in[59]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 6.720 4.000 7.280 ;
    END
  END la_data_in[5]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 201.600 1.000 202.160 4.000 ;
    END
  END la_data_in[60]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 356.160 999.000 356.720 ;
    END
  END la_data_in[61]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 299.040 996.000 299.600 999.000 ;
    END
  END la_data_in[62]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 907.200 996.000 907.760 999.000 ;
    END
  END la_data_in[63]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 870.240 996.000 870.800 999.000 ;
    END
  END la_data_in[6]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 530.880 999.000 531.440 ;
    END
  END la_data_in[7]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 712.320 1.000 712.880 4.000 ;
    END
  END la_data_in[8]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 722.400 4.000 722.960 ;
    END
  END la_data_in[9]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 282.240 996.000 282.800 999.000 ;
    END
  END la_data_out[0]
  PIN la_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 416.640 999.000 417.200 ;
    END
  END la_data_out[10]
  PIN la_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 856.800 4.000 857.360 ;
    END
  END la_data_out[11]
  PIN la_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 551.040 999.000 551.600 ;
    END
  END la_data_out[12]
  PIN la_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 493.920 996.000 494.480 999.000 ;
    END
  END la_data_out[13]
  PIN la_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 443.520 996.000 444.080 999.000 ;
    END
  END la_data_out[14]
  PIN la_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 527.520 1.000 528.080 4.000 ;
    END
  END la_data_out[15]
  PIN la_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 463.680 999.000 464.240 ;
    END
  END la_data_out[16]
  PIN la_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 984.480 996.000 985.040 999.000 ;
    END
  END la_data_out[17]
  PIN la_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 991.200 4.000 991.760 ;
    END
  END la_data_out[18]
  PIN la_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 628.320 999.000 628.880 ;
    END
  END la_data_out[19]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 299.040 1.000 299.600 4.000 ;
    END
  END la_data_out[1]
  PIN la_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 288.960 999.000 289.520 ;
    END
  END la_data_out[20]
  PIN la_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 171.360 4.000 171.920 ;
    END
  END la_data_out[21]
  PIN la_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 127.680 999.000 128.240 ;
    END
  END la_data_out[22]
  PIN la_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 608.160 996.000 608.720 999.000 ;
    END
  END la_data_out[23]
  PIN la_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 792.960 999.000 793.520 ;
    END
  END la_data_out[24]
  PIN la_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 433.440 1.000 434.000 4.000 ;
    END
  END la_data_out[25]
  PIN la_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 779.520 4.000 780.080 ;
    END
  END la_data_out[26]
  PIN la_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 453.600 999.000 454.160 ;
    END
  END la_data_out[27]
  PIN la_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 376.320 4.000 376.880 ;
    END
  END la_data_out[28]
  PIN la_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 588.000 996.000 588.560 999.000 ;
    END
  END la_data_out[29]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 184.800 999.000 185.360 ;
    END
  END la_data_out[2]
  PIN la_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 490.560 1.000 491.120 4.000 ;
    END
  END la_data_out[30]
  PIN la_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 540.960 996.000 541.520 999.000 ;
    END
  END la_data_out[31]
  PIN la_data_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 803.040 999.000 803.600 ;
    END
  END la_data_out[32]
  PIN la_data_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 386.400 999.000 386.960 ;
    END
  END la_data_out[33]
  PIN la_data_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 20.160 999.000 20.720 ;
    END
  END la_data_out[34]
  PIN la_data_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 134.400 999.000 134.960 ;
    END
  END la_data_out[35]
  PIN la_data_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 57.120 4.000 57.680 ;
    END
  END la_data_out[36]
  PIN la_data_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 897.120 4.000 897.680 ;
    END
  END la_data_out[37]
  PIN la_data_out[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 450.240 4.000 450.800 ;
    END
  END la_data_out[38]
  PIN la_data_out[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 840.000 999.000 840.560 ;
    END
  END la_data_out[39]
  PIN la_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 57.120 1.000 57.680 4.000 ;
    END
  END la_data_out[3]
  PIN la_data_out[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 413.280 1.000 413.840 4.000 ;
    END
  END la_data_out[40]
  PIN la_data_out[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 154.560 996.000 155.120 999.000 ;
    END
  END la_data_out[41]
  PIN la_data_out[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 913.920 1.000 914.480 4.000 ;
    END
  END la_data_out[42]
  PIN la_data_out[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 712.320 4.000 712.880 ;
    END
  END la_data_out[43]
  PIN la_data_out[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 228.480 1.000 229.040 4.000 ;
    END
  END la_data_out[44]
  PIN la_data_out[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 903.840 1.000 904.400 4.000 ;
    END
  END la_data_out[45]
  PIN la_data_out[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 571.200 996.000 571.760 999.000 ;
    END
  END la_data_out[46]
  PIN la_data_out[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 349.440 996.000 350.000 999.000 ;
    END
  END la_data_out[47]
  PIN la_data_out[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 964.320 4.000 964.880 ;
    END
  END la_data_out[48]
  PIN la_data_out[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 725.760 996.000 726.320 999.000 ;
    END
  END la_data_out[49]
  PIN la_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 16.800 4.000 17.360 ;
    END
  END la_data_out[4]
  PIN la_data_out[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 782.880 996.000 783.440 999.000 ;
    END
  END la_data_out[50]
  PIN la_data_out[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 426.720 996.000 427.280 999.000 ;
    END
  END la_data_out[51]
  PIN la_data_out[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 144.480 4.000 145.040 ;
    END
  END la_data_out[52]
  PIN la_data_out[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 588.000 999.000 588.560 ;
    END
  END la_data_out[53]
  PIN la_data_out[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 685.440 999.000 686.000 ;
    END
  END la_data_out[54]
  PIN la_data_out[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 887.040 999.000 887.600 ;
    END
  END la_data_out[55]
  PIN la_data_out[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 913.920 4.000 914.480 ;
    END
  END la_data_out[56]
  PIN la_data_out[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 809.760 996.000 810.320 999.000 ;
    END
  END la_data_out[57]
  PIN la_data_out[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 268.800 1.000 269.360 4.000 ;
    END
  END la_data_out[58]
  PIN la_data_out[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 866.880 1.000 867.440 4.000 ;
    END
  END la_data_out[59]
  PIN la_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 67.200 999.000 67.760 ;
    END
  END la_data_out[5]
  PIN la_data_out[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 151.200 4.000 151.760 ;
    END
  END la_data_out[60]
  PIN la_data_out[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 356.160 996.000 356.720 999.000 ;
    END
  END la_data_out[61]
  PIN la_data_out[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 624.960 1.000 625.520 4.000 ;
    END
  END la_data_out[62]
  PIN la_data_out[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 473.760 999.000 474.320 ;
    END
  END la_data_out[63]
  PIN la_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 376.320 999.000 376.880 ;
    END
  END la_data_out[6]
  PIN la_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 705.600 999.000 706.160 ;
    END
  END la_data_out[7]
  PIN la_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 561.120 999.000 561.680 ;
    END
  END la_data_out[8]
  PIN la_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 386.400 996.000 386.960 999.000 ;
    END
  END la_data_out[9]
  PIN la_oenb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 799.680 4.000 800.240 ;
    END
  END la_oenb[0]
  PIN la_oenb[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 732.480 1.000 733.040 4.000 ;
    END
  END la_oenb[10]
  PIN la_oenb[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 876.960 1.000 877.520 4.000 ;
    END
  END la_oenb[11]
  PIN la_oenb[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 144.480 1.000 145.040 4.000 ;
    END
  END la_oenb[12]
  PIN la_oenb[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 124.320 4.000 124.880 ;
    END
  END la_oenb[13]
  PIN la_oenb[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 67.200 996.000 67.760 999.000 ;
    END
  END la_oenb[14]
  PIN la_oenb[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 87.360 999.000 87.920 ;
    END
  END la_oenb[15]
  PIN la_oenb[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 194.880 996.000 195.440 999.000 ;
    END
  END la_oenb[16]
  PIN la_oenb[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 876.960 4.000 877.520 ;
    END
  END la_oenb[17]
  PIN la_oenb[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 880.320 996.000 880.880 999.000 ;
    END
  END la_oenb[18]
  PIN la_oenb[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 742.560 996.000 743.120 999.000 ;
    END
  END la_oenb[19]
  PIN la_oenb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 278.880 1.000 279.440 4.000 ;
    END
  END la_oenb[1]
  PIN la_oenb[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 557.760 4.000 558.320 ;
    END
  END la_oenb[20]
  PIN la_oenb[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 887.040 1.000 887.600 4.000 ;
    END
  END la_oenb[21]
  PIN la_oenb[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 537.600 4.000 538.160 ;
    END
  END la_oenb[22]
  PIN la_oenb[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 181.440 1.000 182.000 4.000 ;
    END
  END la_oenb[23]
  PIN la_oenb[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 614.880 4.000 615.440 ;
    END
  END la_oenb[24]
  PIN la_oenb[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 947.520 999.000 948.080 ;
    END
  END la_oenb[25]
  PIN la_oenb[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 994.560 996.000 995.120 999.000 ;
    END
  END la_oenb[26]
  PIN la_oenb[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 860.160 999.000 860.720 ;
    END
  END la_oenb[27]
  PIN la_oenb[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 819.840 999.000 820.400 ;
    END
  END la_oenb[28]
  PIN la_oenb[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 809.760 999.000 810.320 ;
    END
  END la_oenb[29]
  PIN la_oenb[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 510.720 1.000 511.280 4.000 ;
    END
  END la_oenb[2]
  PIN la_oenb[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 174.720 996.000 175.280 999.000 ;
    END
  END la_oenb[30]
  PIN la_oenb[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 26.880 1.000 27.440 4.000 ;
    END
  END la_oenb[31]
  PIN la_oenb[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 6.720 1.000 7.280 4.000 ;
    END
  END la_oenb[32]
  PIN la_oenb[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 10.080 996.000 10.640 999.000 ;
    END
  END la_oenb[33]
  PIN la_oenb[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 520.800 1.000 521.360 4.000 ;
    END
  END la_oenb[34]
  PIN la_oenb[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 433.440 4.000 434.000 ;
    END
  END la_oenb[35]
  PIN la_oenb[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 547.680 4.000 548.240 ;
    END
  END la_oenb[36]
  PIN la_oenb[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 288.960 4.000 289.520 ;
    END
  END la_oenb[37]
  PIN la_oenb[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 366.240 996.000 366.800 999.000 ;
    END
  END la_oenb[38]
  PIN la_oenb[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 635.040 4.000 635.600 ;
    END
  END la_oenb[39]
  PIN la_oenb[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 191.520 1.000 192.080 4.000 ;
    END
  END la_oenb[3]
  PIN la_oenb[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 443.520 1.000 444.080 4.000 ;
    END
  END la_oenb[40]
  PIN la_oenb[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 500.640 4.000 501.200 ;
    END
  END la_oenb[41]
  PIN la_oenb[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 799.680 1.000 800.240 4.000 ;
    END
  END la_oenb[42]
  PIN la_oenb[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 376.320 1.000 376.880 4.000 ;
    END
  END la_oenb[43]
  PIN la_oenb[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 732.480 4.000 733.040 ;
    END
  END la_oenb[44]
  PIN la_oenb[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 483.840 999.000 484.400 ;
    END
  END la_oenb[45]
  PIN la_oenb[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 665.280 999.000 665.840 ;
    END
  END la_oenb[46]
  PIN la_oenb[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 769.440 1.000 770.000 4.000 ;
    END
  END la_oenb[47]
  PIN la_oenb[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 329.280 996.000 329.840 999.000 ;
    END
  END la_oenb[48]
  PIN la_oenb[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 991.200 1.000 991.760 4.000 ;
    END
  END la_oenb[49]
  PIN la_oenb[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 638.400 999.000 638.960 ;
    END
  END la_oenb[4]
  PIN la_oenb[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 675.360 996.000 675.920 999.000 ;
    END
  END la_oenb[50]
  PIN la_oenb[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 510.720 999.000 511.280 ;
    END
  END la_oenb[51]
  PIN la_oenb[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 759.360 1.000 759.920 4.000 ;
    END
  END la_oenb[52]
  PIN la_oenb[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 887.040 996.000 887.600 999.000 ;
    END
  END la_oenb[53]
  PIN la_oenb[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 97.440 999.000 98.000 ;
    END
  END la_oenb[54]
  PIN la_oenb[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 598.080 996.000 598.640 999.000 ;
    END
  END la_oenb[55]
  PIN la_oenb[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 924.000 1.000 924.560 4.000 ;
    END
  END la_oenb[56]
  PIN la_oenb[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 490.560 4.000 491.120 ;
    END
  END la_oenb[57]
  PIN la_oenb[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 124.320 1.000 124.880 4.000 ;
    END
  END la_oenb[58]
  PIN la_oenb[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 504.000 999.000 504.560 ;
    END
  END la_oenb[59]
  PIN la_oenb[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 954.240 4.000 954.800 ;
    END
  END la_oenb[5]
  PIN la_oenb[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 658.560 999.000 659.120 ;
    END
  END la_oenb[60]
  PIN la_oenb[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 248.640 1.000 249.200 4.000 ;
    END
  END la_oenb[61]
  PIN la_oenb[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 954.240 1.000 954.800 4.000 ;
    END
  END la_oenb[62]
  PIN la_oenb[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 181.440 4.000 182.000 ;
    END
  END la_oenb[63]
  PIN la_oenb[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 860.160 996.000 860.720 999.000 ;
    END
  END la_oenb[6]
  PIN la_oenb[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 762.720 999.000 763.280 ;
    END
  END la_oenb[7]
  PIN la_oenb[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 252.000 996.000 252.560 999.000 ;
    END
  END la_oenb[8]
  PIN la_oenb[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 645.120 4.000 645.680 ;
    END
  END la_oenb[9]
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 22.240 15.380 23.840 984.220 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 175.840 15.380 177.440 984.220 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 329.440 15.380 331.040 984.220 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 483.040 15.380 484.640 984.220 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 636.640 15.380 638.240 984.220 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 790.240 15.380 791.840 984.220 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 943.840 15.380 945.440 984.220 ;
    END
  END vdd
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 99.040 15.380 100.640 984.220 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 252.640 15.380 254.240 984.220 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 406.240 15.380 407.840 984.220 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 559.840 15.380 561.440 984.220 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 713.440 15.380 715.040 984.220 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 867.040 15.380 868.640 984.220 ;
    END
  END vss
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 174.720 999.000 175.280 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 184.800 996.000 185.360 999.000 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 349.440 999.000 350.000 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 665.280 996.000 665.840 999.000 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 453.600 996.000 454.160 999.000 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 57.120 996.000 57.680 999.000 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 84.000 1.000 84.560 4.000 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 557.760 1.000 558.320 4.000 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 735.840 999.000 736.400 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 675.360 999.000 675.920 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 635.040 1.000 635.600 4.000 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 598.080 999.000 598.640 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 309.120 999.000 309.680 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 964.320 1.000 964.880 4.000 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 67.200 4.000 67.760 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 588.000 4.000 588.560 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 567.840 1.000 568.400 4.000 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 809.760 1.000 810.320 4.000 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 231.840 999.000 232.400 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 117.600 996.000 118.160 999.000 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 547.680 1.000 548.240 4.000 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 104.160 1.000 104.720 4.000 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 339.360 996.000 339.920 999.000 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 581.280 999.000 581.840 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 957.600 999.000 958.160 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 114.240 4.000 114.800 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 393.120 4.000 393.680 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 426.720 999.000 427.280 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 779.520 1.000 780.080 4.000 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 772.800 996.000 773.360 999.000 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 752.640 1.000 753.200 4.000 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 480.480 4.000 481.040 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 47.040 1.000 47.600 4.000 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 0.000 999.000 0.560 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 272.160 999.000 272.720 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 319.200 996.000 319.760 999.000 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 870.240 999.000 870.800 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 769.440 4.000 770.000 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 846.720 4.000 847.280 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 809.760 4.000 810.320 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 36.960 1.000 37.520 4.000 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 211.680 4.000 212.240 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 520.800 999.000 521.360 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 577.920 1.000 578.480 4.000 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 685.440 996.000 686.000 999.000 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 927.360 996.000 927.920 999.000 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 50.400 996.000 50.960 999.000 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 151.200 1.000 151.760 4.000 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 248.640 4.000 249.200 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 957.600 996.000 958.160 999.000 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 598.080 4.000 598.640 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 782.880 999.000 783.440 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 329.280 999.000 329.840 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 692.160 1.000 692.720 4.000 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 829.920 996.000 830.480 999.000 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 241.920 996.000 242.480 999.000 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 315.840 1.000 316.400 4.000 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 608.160 999.000 608.720 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 819.840 1.000 820.400 4.000 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 299.040 999.000 299.600 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 527.520 4.000 528.080 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 40.320 999.000 40.880 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 161.280 1.000 161.840 4.000 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 500.640 1.000 501.200 4.000 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 433.440 999.000 434.000 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 792.960 996.000 793.520 999.000 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 897.120 999.000 897.680 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 50.400 999.000 50.960 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 201.600 4.000 202.160 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 571.200 999.000 571.760 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 16.800 1.000 17.360 4.000 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 917.280 999.000 917.840 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 752.640 996.000 753.200 999.000 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 117.600 999.000 118.160 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 715.680 996.000 716.240 999.000 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 278.880 4.000 279.440 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 315.840 4.000 316.400 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 675.360 1.000 675.920 4.000 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 0.000 1.000 0.560 4.000 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 789.600 1.000 790.160 4.000 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 470.400 4.000 470.960 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 866.880 4.000 867.440 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 272.160 996.000 272.720 999.000 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 325.920 4.000 326.480 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 211.680 1.000 212.240 4.000 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 73.920 1.000 74.480 4.000 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 520.800 996.000 521.360 999.000 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 288.960 996.000 289.520 999.000 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 537.600 1.000 538.160 4.000 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 695.520 996.000 696.080 999.000 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 282.240 999.000 282.800 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 655.200 4.000 655.760 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 772.800 999.000 773.360 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 221.760 1.000 222.320 4.000 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 383.040 1.000 383.600 4.000 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 84.000 4.000 84.560 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 742.560 999.000 743.120 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 604.800 1.000 605.360 4.000 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 658.560 996.000 659.120 999.000 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 648.480 996.000 649.040 999.000 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 924.000 4.000 924.560 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 107.520 996.000 108.080 999.000 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 722.400 1.000 722.960 4.000 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 221.760 4.000 222.320 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 1.000 829.920 4.000 830.480 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 996.000 493.920 999.000 494.480 ;
    END
  END wbs_we_i
  OBS
      LAYER Metal1 ;
        RECT 6.720 8.550 992.880 984.220 ;
      LAYER Metal2 ;
        RECT 0.860 995.700 9.780 996.660 ;
        RECT 10.940 995.700 19.860 996.660 ;
        RECT 21.020 995.700 29.940 996.660 ;
        RECT 31.100 995.700 40.020 996.660 ;
        RECT 41.180 995.700 50.100 996.660 ;
        RECT 51.260 995.700 56.820 996.660 ;
        RECT 57.980 995.700 66.900 996.660 ;
        RECT 68.060 995.700 76.980 996.660 ;
        RECT 78.140 995.700 87.060 996.660 ;
        RECT 88.220 995.700 97.140 996.660 ;
        RECT 98.300 995.700 107.220 996.660 ;
        RECT 108.380 995.700 117.300 996.660 ;
        RECT 118.460 995.700 127.380 996.660 ;
        RECT 128.540 995.700 134.100 996.660 ;
        RECT 135.260 995.700 144.180 996.660 ;
        RECT 145.340 995.700 154.260 996.660 ;
        RECT 155.420 995.700 164.340 996.660 ;
        RECT 165.500 995.700 174.420 996.660 ;
        RECT 175.580 995.700 184.500 996.660 ;
        RECT 185.660 995.700 194.580 996.660 ;
        RECT 195.740 995.700 204.660 996.660 ;
        RECT 205.820 995.700 211.380 996.660 ;
        RECT 212.540 995.700 221.460 996.660 ;
        RECT 222.620 995.700 231.540 996.660 ;
        RECT 232.700 995.700 241.620 996.660 ;
        RECT 242.780 995.700 251.700 996.660 ;
        RECT 252.860 995.700 261.780 996.660 ;
        RECT 262.940 995.700 271.860 996.660 ;
        RECT 273.020 995.700 281.940 996.660 ;
        RECT 283.100 995.700 288.660 996.660 ;
        RECT 289.820 995.700 298.740 996.660 ;
        RECT 299.900 995.700 308.820 996.660 ;
        RECT 309.980 995.700 318.900 996.660 ;
        RECT 320.060 995.700 328.980 996.660 ;
        RECT 330.140 995.700 339.060 996.660 ;
        RECT 340.220 995.700 349.140 996.660 ;
        RECT 350.300 995.700 355.860 996.660 ;
        RECT 357.020 995.700 365.940 996.660 ;
        RECT 367.100 995.700 376.020 996.660 ;
        RECT 377.180 995.700 386.100 996.660 ;
        RECT 387.260 995.700 396.180 996.660 ;
        RECT 397.340 995.700 406.260 996.660 ;
        RECT 407.420 995.700 416.340 996.660 ;
        RECT 417.500 995.700 426.420 996.660 ;
        RECT 427.580 995.700 433.140 996.660 ;
        RECT 434.300 995.700 443.220 996.660 ;
        RECT 444.380 995.700 453.300 996.660 ;
        RECT 454.460 995.700 463.380 996.660 ;
        RECT 464.540 995.700 473.460 996.660 ;
        RECT 474.620 995.700 483.540 996.660 ;
        RECT 484.700 995.700 493.620 996.660 ;
        RECT 494.780 995.700 503.700 996.660 ;
        RECT 504.860 995.700 510.420 996.660 ;
        RECT 511.580 995.700 520.500 996.660 ;
        RECT 521.660 995.700 530.580 996.660 ;
        RECT 531.740 995.700 540.660 996.660 ;
        RECT 541.820 995.700 550.740 996.660 ;
        RECT 551.900 995.700 560.820 996.660 ;
        RECT 561.980 995.700 570.900 996.660 ;
        RECT 572.060 995.700 580.980 996.660 ;
        RECT 582.140 995.700 587.700 996.660 ;
        RECT 588.860 995.700 597.780 996.660 ;
        RECT 598.940 995.700 607.860 996.660 ;
        RECT 609.020 995.700 617.940 996.660 ;
        RECT 619.100 995.700 628.020 996.660 ;
        RECT 629.180 995.700 638.100 996.660 ;
        RECT 639.260 995.700 648.180 996.660 ;
        RECT 649.340 995.700 658.260 996.660 ;
        RECT 659.420 995.700 664.980 996.660 ;
        RECT 666.140 995.700 675.060 996.660 ;
        RECT 676.220 995.700 685.140 996.660 ;
        RECT 686.300 995.700 695.220 996.660 ;
        RECT 696.380 995.700 705.300 996.660 ;
        RECT 706.460 995.700 715.380 996.660 ;
        RECT 716.540 995.700 725.460 996.660 ;
        RECT 726.620 995.700 735.540 996.660 ;
        RECT 736.700 995.700 742.260 996.660 ;
        RECT 743.420 995.700 752.340 996.660 ;
        RECT 753.500 995.700 762.420 996.660 ;
        RECT 763.580 995.700 772.500 996.660 ;
        RECT 773.660 995.700 782.580 996.660 ;
        RECT 783.740 995.700 792.660 996.660 ;
        RECT 793.820 995.700 802.740 996.660 ;
        RECT 803.900 995.700 809.460 996.660 ;
        RECT 810.620 995.700 819.540 996.660 ;
        RECT 820.700 995.700 829.620 996.660 ;
        RECT 830.780 995.700 839.700 996.660 ;
        RECT 840.860 995.700 849.780 996.660 ;
        RECT 850.940 995.700 859.860 996.660 ;
        RECT 861.020 995.700 869.940 996.660 ;
        RECT 871.100 995.700 880.020 996.660 ;
        RECT 881.180 995.700 886.740 996.660 ;
        RECT 887.900 995.700 896.820 996.660 ;
        RECT 897.980 995.700 906.900 996.660 ;
        RECT 908.060 995.700 916.980 996.660 ;
        RECT 918.140 995.700 927.060 996.660 ;
        RECT 928.220 995.700 937.140 996.660 ;
        RECT 938.300 995.700 947.220 996.660 ;
        RECT 948.380 995.700 957.300 996.660 ;
        RECT 958.460 995.700 964.020 996.660 ;
        RECT 965.180 995.700 974.100 996.660 ;
        RECT 975.260 995.700 984.180 996.660 ;
        RECT 985.340 995.700 990.500 996.660 ;
        RECT 0.140 4.300 990.500 995.700 ;
        RECT 0.860 4.000 6.420 4.300 ;
        RECT 7.580 4.000 16.500 4.300 ;
        RECT 17.660 4.000 26.580 4.300 ;
        RECT 27.740 4.000 36.660 4.300 ;
        RECT 37.820 4.000 46.740 4.300 ;
        RECT 47.900 4.000 56.820 4.300 ;
        RECT 57.980 4.000 66.900 4.300 ;
        RECT 68.060 4.000 73.620 4.300 ;
        RECT 74.780 4.000 83.700 4.300 ;
        RECT 84.860 4.000 93.780 4.300 ;
        RECT 94.940 4.000 103.860 4.300 ;
        RECT 105.020 4.000 113.940 4.300 ;
        RECT 115.100 4.000 124.020 4.300 ;
        RECT 125.180 4.000 134.100 4.300 ;
        RECT 135.260 4.000 144.180 4.300 ;
        RECT 145.340 4.000 150.900 4.300 ;
        RECT 152.060 4.000 160.980 4.300 ;
        RECT 162.140 4.000 171.060 4.300 ;
        RECT 172.220 4.000 181.140 4.300 ;
        RECT 182.300 4.000 191.220 4.300 ;
        RECT 192.380 4.000 201.300 4.300 ;
        RECT 202.460 4.000 211.380 4.300 ;
        RECT 212.540 4.000 221.460 4.300 ;
        RECT 222.620 4.000 228.180 4.300 ;
        RECT 229.340 4.000 238.260 4.300 ;
        RECT 239.420 4.000 248.340 4.300 ;
        RECT 249.500 4.000 258.420 4.300 ;
        RECT 259.580 4.000 268.500 4.300 ;
        RECT 269.660 4.000 278.580 4.300 ;
        RECT 279.740 4.000 288.660 4.300 ;
        RECT 289.820 4.000 298.740 4.300 ;
        RECT 299.900 4.000 305.460 4.300 ;
        RECT 306.620 4.000 315.540 4.300 ;
        RECT 316.700 4.000 325.620 4.300 ;
        RECT 326.780 4.000 335.700 4.300 ;
        RECT 336.860 4.000 345.780 4.300 ;
        RECT 346.940 4.000 355.860 4.300 ;
        RECT 357.020 4.000 365.940 4.300 ;
        RECT 367.100 4.000 376.020 4.300 ;
        RECT 377.180 4.000 382.740 4.300 ;
        RECT 383.900 4.000 392.820 4.300 ;
        RECT 393.980 4.000 402.900 4.300 ;
        RECT 404.060 4.000 412.980 4.300 ;
        RECT 414.140 4.000 423.060 4.300 ;
        RECT 424.220 4.000 433.140 4.300 ;
        RECT 434.300 4.000 443.220 4.300 ;
        RECT 444.380 4.000 449.940 4.300 ;
        RECT 451.100 4.000 460.020 4.300 ;
        RECT 461.180 4.000 470.100 4.300 ;
        RECT 471.260 4.000 480.180 4.300 ;
        RECT 481.340 4.000 490.260 4.300 ;
        RECT 491.420 4.000 500.340 4.300 ;
        RECT 501.500 4.000 510.420 4.300 ;
        RECT 511.580 4.000 520.500 4.300 ;
        RECT 521.660 4.000 527.220 4.300 ;
        RECT 528.380 4.000 537.300 4.300 ;
        RECT 538.460 4.000 547.380 4.300 ;
        RECT 548.540 4.000 557.460 4.300 ;
        RECT 558.620 4.000 567.540 4.300 ;
        RECT 568.700 4.000 577.620 4.300 ;
        RECT 578.780 4.000 587.700 4.300 ;
        RECT 588.860 4.000 597.780 4.300 ;
        RECT 598.940 4.000 604.500 4.300 ;
        RECT 605.660 4.000 614.580 4.300 ;
        RECT 615.740 4.000 624.660 4.300 ;
        RECT 625.820 4.000 634.740 4.300 ;
        RECT 635.900 4.000 644.820 4.300 ;
        RECT 645.980 4.000 654.900 4.300 ;
        RECT 656.060 4.000 664.980 4.300 ;
        RECT 666.140 4.000 675.060 4.300 ;
        RECT 676.220 4.000 681.780 4.300 ;
        RECT 682.940 4.000 691.860 4.300 ;
        RECT 693.020 4.000 701.940 4.300 ;
        RECT 703.100 4.000 712.020 4.300 ;
        RECT 713.180 4.000 722.100 4.300 ;
        RECT 723.260 4.000 732.180 4.300 ;
        RECT 733.340 4.000 742.260 4.300 ;
        RECT 743.420 4.000 752.340 4.300 ;
        RECT 753.500 4.000 759.060 4.300 ;
        RECT 760.220 4.000 769.140 4.300 ;
        RECT 770.300 4.000 779.220 4.300 ;
        RECT 780.380 4.000 789.300 4.300 ;
        RECT 790.460 4.000 799.380 4.300 ;
        RECT 800.540 4.000 809.460 4.300 ;
        RECT 810.620 4.000 819.540 4.300 ;
        RECT 820.700 4.000 829.620 4.300 ;
        RECT 830.780 4.000 836.340 4.300 ;
        RECT 837.500 4.000 846.420 4.300 ;
        RECT 847.580 4.000 856.500 4.300 ;
        RECT 857.660 4.000 866.580 4.300 ;
        RECT 867.740 4.000 876.660 4.300 ;
        RECT 877.820 4.000 886.740 4.300 ;
        RECT 887.900 4.000 896.820 4.300 ;
        RECT 897.980 4.000 903.540 4.300 ;
        RECT 904.700 4.000 913.620 4.300 ;
        RECT 914.780 4.000 923.700 4.300 ;
        RECT 924.860 4.000 933.780 4.300 ;
        RECT 934.940 4.000 943.860 4.300 ;
        RECT 945.020 4.000 953.940 4.300 ;
        RECT 955.100 4.000 964.020 4.300 ;
        RECT 965.180 4.000 974.100 4.300 ;
        RECT 975.260 4.000 980.820 4.300 ;
        RECT 981.980 4.000 990.500 4.300 ;
      LAYER Metal3 ;
        RECT 0.090 994.260 995.700 994.980 ;
        RECT 0.090 992.060 996.660 994.260 ;
        RECT 0.090 990.900 0.700 992.060 ;
        RECT 4.300 990.900 996.660 992.060 ;
        RECT 0.090 985.340 996.660 990.900 ;
        RECT 0.090 984.180 995.700 985.340 ;
        RECT 0.090 981.980 996.660 984.180 ;
        RECT 0.090 980.820 0.700 981.980 ;
        RECT 4.300 980.820 996.660 981.980 ;
        RECT 0.090 975.260 996.660 980.820 ;
        RECT 0.090 974.100 0.700 975.260 ;
        RECT 4.300 974.100 995.700 975.260 ;
        RECT 0.090 965.180 996.660 974.100 ;
        RECT 0.090 964.020 0.700 965.180 ;
        RECT 4.300 964.020 995.700 965.180 ;
        RECT 0.090 958.460 996.660 964.020 ;
        RECT 0.090 957.300 995.700 958.460 ;
        RECT 0.090 955.100 996.660 957.300 ;
        RECT 0.090 953.940 0.700 955.100 ;
        RECT 4.300 953.940 996.660 955.100 ;
        RECT 0.090 948.380 996.660 953.940 ;
        RECT 0.090 947.220 995.700 948.380 ;
        RECT 0.090 945.020 996.660 947.220 ;
        RECT 0.090 943.860 0.700 945.020 ;
        RECT 4.300 943.860 996.660 945.020 ;
        RECT 0.090 938.300 996.660 943.860 ;
        RECT 0.090 937.140 995.700 938.300 ;
        RECT 0.090 934.940 996.660 937.140 ;
        RECT 0.090 933.780 0.700 934.940 ;
        RECT 4.300 933.780 996.660 934.940 ;
        RECT 0.090 928.220 996.660 933.780 ;
        RECT 0.090 927.060 995.700 928.220 ;
        RECT 0.090 924.860 996.660 927.060 ;
        RECT 0.090 923.700 0.700 924.860 ;
        RECT 4.300 923.700 996.660 924.860 ;
        RECT 0.090 918.140 996.660 923.700 ;
        RECT 0.090 916.980 995.700 918.140 ;
        RECT 0.090 914.780 996.660 916.980 ;
        RECT 0.090 913.620 0.700 914.780 ;
        RECT 4.300 913.620 996.660 914.780 ;
        RECT 0.090 908.060 996.660 913.620 ;
        RECT 0.090 906.900 995.700 908.060 ;
        RECT 0.090 904.700 996.660 906.900 ;
        RECT 0.090 903.540 0.700 904.700 ;
        RECT 4.300 903.540 996.660 904.700 ;
        RECT 0.090 897.980 996.660 903.540 ;
        RECT 0.090 896.820 0.700 897.980 ;
        RECT 4.300 896.820 995.700 897.980 ;
        RECT 0.090 887.900 996.660 896.820 ;
        RECT 0.090 886.740 0.700 887.900 ;
        RECT 4.300 886.740 995.700 887.900 ;
        RECT 0.090 881.180 996.660 886.740 ;
        RECT 0.090 880.020 995.700 881.180 ;
        RECT 0.090 877.820 996.660 880.020 ;
        RECT 0.090 876.660 0.700 877.820 ;
        RECT 4.300 876.660 996.660 877.820 ;
        RECT 0.090 871.100 996.660 876.660 ;
        RECT 0.090 869.940 995.700 871.100 ;
        RECT 0.090 867.740 996.660 869.940 ;
        RECT 0.090 866.580 0.700 867.740 ;
        RECT 4.300 866.580 996.660 867.740 ;
        RECT 0.090 861.020 996.660 866.580 ;
        RECT 0.090 859.860 995.700 861.020 ;
        RECT 0.090 857.660 996.660 859.860 ;
        RECT 0.090 856.500 0.700 857.660 ;
        RECT 4.300 856.500 996.660 857.660 ;
        RECT 0.090 850.940 996.660 856.500 ;
        RECT 0.090 849.780 995.700 850.940 ;
        RECT 0.090 847.580 996.660 849.780 ;
        RECT 0.090 846.420 0.700 847.580 ;
        RECT 4.300 846.420 996.660 847.580 ;
        RECT 0.090 840.860 996.660 846.420 ;
        RECT 0.090 839.700 995.700 840.860 ;
        RECT 0.090 837.500 996.660 839.700 ;
        RECT 0.090 836.340 0.700 837.500 ;
        RECT 4.300 836.340 996.660 837.500 ;
        RECT 0.090 830.780 996.660 836.340 ;
        RECT 0.090 829.620 0.700 830.780 ;
        RECT 4.300 829.620 995.700 830.780 ;
        RECT 0.090 820.700 996.660 829.620 ;
        RECT 0.090 819.540 0.700 820.700 ;
        RECT 4.300 819.540 995.700 820.700 ;
        RECT 0.090 810.620 996.660 819.540 ;
        RECT 0.090 809.460 0.700 810.620 ;
        RECT 4.300 809.460 995.700 810.620 ;
        RECT 0.090 803.900 996.660 809.460 ;
        RECT 0.090 802.740 995.700 803.900 ;
        RECT 0.090 800.540 996.660 802.740 ;
        RECT 0.090 799.380 0.700 800.540 ;
        RECT 4.300 799.380 996.660 800.540 ;
        RECT 0.090 793.820 996.660 799.380 ;
        RECT 0.090 792.660 995.700 793.820 ;
        RECT 0.090 790.460 996.660 792.660 ;
        RECT 0.090 789.300 0.700 790.460 ;
        RECT 4.300 789.300 996.660 790.460 ;
        RECT 0.090 783.740 996.660 789.300 ;
        RECT 0.090 782.580 995.700 783.740 ;
        RECT 0.090 780.380 996.660 782.580 ;
        RECT 0.090 779.220 0.700 780.380 ;
        RECT 4.300 779.220 996.660 780.380 ;
        RECT 0.090 773.660 996.660 779.220 ;
        RECT 0.090 772.500 995.700 773.660 ;
        RECT 0.090 770.300 996.660 772.500 ;
        RECT 0.090 769.140 0.700 770.300 ;
        RECT 4.300 769.140 996.660 770.300 ;
        RECT 0.090 763.580 996.660 769.140 ;
        RECT 0.090 762.420 995.700 763.580 ;
        RECT 0.090 760.220 996.660 762.420 ;
        RECT 0.090 759.060 0.700 760.220 ;
        RECT 4.300 759.060 996.660 760.220 ;
        RECT 0.090 753.500 996.660 759.060 ;
        RECT 0.090 752.340 0.700 753.500 ;
        RECT 4.300 752.340 995.700 753.500 ;
        RECT 0.090 743.420 996.660 752.340 ;
        RECT 0.090 742.260 0.700 743.420 ;
        RECT 4.300 742.260 995.700 743.420 ;
        RECT 0.090 736.700 996.660 742.260 ;
        RECT 0.090 735.540 995.700 736.700 ;
        RECT 0.090 733.340 996.660 735.540 ;
        RECT 0.090 732.180 0.700 733.340 ;
        RECT 4.300 732.180 996.660 733.340 ;
        RECT 0.090 726.620 996.660 732.180 ;
        RECT 0.090 725.460 995.700 726.620 ;
        RECT 0.090 723.260 996.660 725.460 ;
        RECT 0.090 722.100 0.700 723.260 ;
        RECT 4.300 722.100 996.660 723.260 ;
        RECT 0.090 716.540 996.660 722.100 ;
        RECT 0.090 715.380 995.700 716.540 ;
        RECT 0.090 713.180 996.660 715.380 ;
        RECT 0.090 712.020 0.700 713.180 ;
        RECT 4.300 712.020 996.660 713.180 ;
        RECT 0.090 706.460 996.660 712.020 ;
        RECT 0.090 705.300 995.700 706.460 ;
        RECT 0.090 703.100 996.660 705.300 ;
        RECT 0.090 701.940 0.700 703.100 ;
        RECT 4.300 701.940 996.660 703.100 ;
        RECT 0.090 696.380 996.660 701.940 ;
        RECT 0.090 695.220 995.700 696.380 ;
        RECT 0.090 693.020 996.660 695.220 ;
        RECT 0.090 691.860 0.700 693.020 ;
        RECT 4.300 691.860 996.660 693.020 ;
        RECT 0.090 686.300 996.660 691.860 ;
        RECT 0.090 685.140 995.700 686.300 ;
        RECT 0.090 682.940 996.660 685.140 ;
        RECT 0.090 681.780 0.700 682.940 ;
        RECT 4.300 681.780 996.660 682.940 ;
        RECT 0.090 676.220 996.660 681.780 ;
        RECT 0.090 675.060 0.700 676.220 ;
        RECT 4.300 675.060 995.700 676.220 ;
        RECT 0.090 666.140 996.660 675.060 ;
        RECT 0.090 664.980 0.700 666.140 ;
        RECT 4.300 664.980 995.700 666.140 ;
        RECT 0.090 659.420 996.660 664.980 ;
        RECT 0.090 658.260 995.700 659.420 ;
        RECT 0.090 656.060 996.660 658.260 ;
        RECT 0.090 654.900 0.700 656.060 ;
        RECT 4.300 654.900 996.660 656.060 ;
        RECT 0.090 649.340 996.660 654.900 ;
        RECT 0.090 648.180 995.700 649.340 ;
        RECT 0.090 645.980 996.660 648.180 ;
        RECT 0.090 644.820 0.700 645.980 ;
        RECT 4.300 644.820 996.660 645.980 ;
        RECT 0.090 639.260 996.660 644.820 ;
        RECT 0.090 638.100 995.700 639.260 ;
        RECT 0.090 635.900 996.660 638.100 ;
        RECT 0.090 634.740 0.700 635.900 ;
        RECT 4.300 634.740 996.660 635.900 ;
        RECT 0.090 629.180 996.660 634.740 ;
        RECT 0.090 628.020 995.700 629.180 ;
        RECT 0.090 625.820 996.660 628.020 ;
        RECT 0.090 624.660 0.700 625.820 ;
        RECT 4.300 624.660 996.660 625.820 ;
        RECT 0.090 619.100 996.660 624.660 ;
        RECT 0.090 617.940 995.700 619.100 ;
        RECT 0.090 615.740 996.660 617.940 ;
        RECT 0.090 614.580 0.700 615.740 ;
        RECT 4.300 614.580 996.660 615.740 ;
        RECT 0.090 609.020 996.660 614.580 ;
        RECT 0.090 607.860 995.700 609.020 ;
        RECT 0.090 605.660 996.660 607.860 ;
        RECT 0.090 604.500 0.700 605.660 ;
        RECT 4.300 604.500 996.660 605.660 ;
        RECT 0.090 598.940 996.660 604.500 ;
        RECT 0.090 597.780 0.700 598.940 ;
        RECT 4.300 597.780 995.700 598.940 ;
        RECT 0.090 588.860 996.660 597.780 ;
        RECT 0.090 587.700 0.700 588.860 ;
        RECT 4.300 587.700 995.700 588.860 ;
        RECT 0.090 582.140 996.660 587.700 ;
        RECT 0.090 580.980 995.700 582.140 ;
        RECT 0.090 578.780 996.660 580.980 ;
        RECT 0.090 577.620 0.700 578.780 ;
        RECT 4.300 577.620 996.660 578.780 ;
        RECT 0.090 572.060 996.660 577.620 ;
        RECT 0.090 570.900 995.700 572.060 ;
        RECT 0.090 568.700 996.660 570.900 ;
        RECT 0.090 567.540 0.700 568.700 ;
        RECT 4.300 567.540 996.660 568.700 ;
        RECT 0.090 561.980 996.660 567.540 ;
        RECT 0.090 560.820 995.700 561.980 ;
        RECT 0.090 558.620 996.660 560.820 ;
        RECT 0.090 557.460 0.700 558.620 ;
        RECT 4.300 557.460 996.660 558.620 ;
        RECT 0.090 551.900 996.660 557.460 ;
        RECT 0.090 550.740 995.700 551.900 ;
        RECT 0.090 548.540 996.660 550.740 ;
        RECT 0.090 547.380 0.700 548.540 ;
        RECT 4.300 547.380 996.660 548.540 ;
        RECT 0.090 541.820 996.660 547.380 ;
        RECT 0.090 540.660 995.700 541.820 ;
        RECT 0.090 538.460 996.660 540.660 ;
        RECT 0.090 537.300 0.700 538.460 ;
        RECT 4.300 537.300 996.660 538.460 ;
        RECT 0.090 531.740 996.660 537.300 ;
        RECT 0.090 530.580 995.700 531.740 ;
        RECT 0.090 528.380 996.660 530.580 ;
        RECT 0.090 527.220 0.700 528.380 ;
        RECT 4.300 527.220 996.660 528.380 ;
        RECT 0.090 521.660 996.660 527.220 ;
        RECT 0.090 520.500 0.700 521.660 ;
        RECT 4.300 520.500 995.700 521.660 ;
        RECT 0.090 511.580 996.660 520.500 ;
        RECT 0.090 510.420 0.700 511.580 ;
        RECT 4.300 510.420 995.700 511.580 ;
        RECT 0.090 504.860 996.660 510.420 ;
        RECT 0.090 503.700 995.700 504.860 ;
        RECT 0.090 501.500 996.660 503.700 ;
        RECT 0.090 500.340 0.700 501.500 ;
        RECT 4.300 500.340 996.660 501.500 ;
        RECT 0.090 494.780 996.660 500.340 ;
        RECT 0.090 493.620 995.700 494.780 ;
        RECT 0.090 491.420 996.660 493.620 ;
        RECT 0.090 490.260 0.700 491.420 ;
        RECT 4.300 490.260 996.660 491.420 ;
        RECT 0.090 484.700 996.660 490.260 ;
        RECT 0.090 483.540 995.700 484.700 ;
        RECT 0.090 481.340 996.660 483.540 ;
        RECT 0.090 480.180 0.700 481.340 ;
        RECT 4.300 480.180 996.660 481.340 ;
        RECT 0.090 474.620 996.660 480.180 ;
        RECT 0.090 473.460 995.700 474.620 ;
        RECT 0.090 471.260 996.660 473.460 ;
        RECT 0.090 470.100 0.700 471.260 ;
        RECT 4.300 470.100 996.660 471.260 ;
        RECT 0.090 464.540 996.660 470.100 ;
        RECT 0.090 463.380 995.700 464.540 ;
        RECT 0.090 461.180 996.660 463.380 ;
        RECT 0.090 460.020 0.700 461.180 ;
        RECT 4.300 460.020 996.660 461.180 ;
        RECT 0.090 454.460 996.660 460.020 ;
        RECT 0.090 453.300 995.700 454.460 ;
        RECT 0.090 451.100 996.660 453.300 ;
        RECT 0.090 449.940 0.700 451.100 ;
        RECT 4.300 449.940 996.660 451.100 ;
        RECT 0.090 444.380 996.660 449.940 ;
        RECT 0.090 443.220 0.700 444.380 ;
        RECT 4.300 443.220 995.700 444.380 ;
        RECT 0.090 434.300 996.660 443.220 ;
        RECT 0.090 433.140 0.700 434.300 ;
        RECT 4.300 433.140 995.700 434.300 ;
        RECT 0.090 427.580 996.660 433.140 ;
        RECT 0.090 426.420 995.700 427.580 ;
        RECT 0.090 424.220 996.660 426.420 ;
        RECT 0.090 423.060 0.700 424.220 ;
        RECT 4.300 423.060 996.660 424.220 ;
        RECT 0.090 417.500 996.660 423.060 ;
        RECT 0.090 416.340 995.700 417.500 ;
        RECT 0.090 414.140 996.660 416.340 ;
        RECT 0.090 412.980 0.700 414.140 ;
        RECT 4.300 412.980 996.660 414.140 ;
        RECT 0.090 407.420 996.660 412.980 ;
        RECT 0.090 406.260 995.700 407.420 ;
        RECT 0.090 404.060 996.660 406.260 ;
        RECT 0.090 402.900 0.700 404.060 ;
        RECT 4.300 402.900 996.660 404.060 ;
        RECT 0.090 397.340 996.660 402.900 ;
        RECT 0.090 396.180 995.700 397.340 ;
        RECT 0.090 393.980 996.660 396.180 ;
        RECT 0.090 392.820 0.700 393.980 ;
        RECT 4.300 392.820 996.660 393.980 ;
        RECT 0.090 387.260 996.660 392.820 ;
        RECT 0.090 386.100 995.700 387.260 ;
        RECT 0.090 383.900 996.660 386.100 ;
        RECT 0.090 382.740 0.700 383.900 ;
        RECT 4.300 382.740 996.660 383.900 ;
        RECT 0.090 377.180 996.660 382.740 ;
        RECT 0.090 376.020 0.700 377.180 ;
        RECT 4.300 376.020 995.700 377.180 ;
        RECT 0.090 367.100 996.660 376.020 ;
        RECT 0.090 365.940 0.700 367.100 ;
        RECT 4.300 365.940 995.700 367.100 ;
        RECT 0.090 357.020 996.660 365.940 ;
        RECT 0.090 355.860 0.700 357.020 ;
        RECT 4.300 355.860 995.700 357.020 ;
        RECT 0.090 350.300 996.660 355.860 ;
        RECT 0.090 349.140 995.700 350.300 ;
        RECT 0.090 346.940 996.660 349.140 ;
        RECT 0.090 345.780 0.700 346.940 ;
        RECT 4.300 345.780 996.660 346.940 ;
        RECT 0.090 340.220 996.660 345.780 ;
        RECT 0.090 339.060 995.700 340.220 ;
        RECT 0.090 336.860 996.660 339.060 ;
        RECT 0.090 335.700 0.700 336.860 ;
        RECT 4.300 335.700 996.660 336.860 ;
        RECT 0.090 330.140 996.660 335.700 ;
        RECT 0.090 328.980 995.700 330.140 ;
        RECT 0.090 326.780 996.660 328.980 ;
        RECT 0.090 325.620 0.700 326.780 ;
        RECT 4.300 325.620 996.660 326.780 ;
        RECT 0.090 320.060 996.660 325.620 ;
        RECT 0.090 318.900 995.700 320.060 ;
        RECT 0.090 316.700 996.660 318.900 ;
        RECT 0.090 315.540 0.700 316.700 ;
        RECT 4.300 315.540 996.660 316.700 ;
        RECT 0.090 309.980 996.660 315.540 ;
        RECT 0.090 308.820 995.700 309.980 ;
        RECT 0.090 306.620 996.660 308.820 ;
        RECT 0.090 305.460 0.700 306.620 ;
        RECT 4.300 305.460 996.660 306.620 ;
        RECT 0.090 299.900 996.660 305.460 ;
        RECT 0.090 298.740 0.700 299.900 ;
        RECT 4.300 298.740 995.700 299.900 ;
        RECT 0.090 289.820 996.660 298.740 ;
        RECT 0.090 288.660 0.700 289.820 ;
        RECT 4.300 288.660 995.700 289.820 ;
        RECT 0.090 283.100 996.660 288.660 ;
        RECT 0.090 281.940 995.700 283.100 ;
        RECT 0.090 279.740 996.660 281.940 ;
        RECT 0.090 278.580 0.700 279.740 ;
        RECT 4.300 278.580 996.660 279.740 ;
        RECT 0.090 273.020 996.660 278.580 ;
        RECT 0.090 271.860 995.700 273.020 ;
        RECT 0.090 269.660 996.660 271.860 ;
        RECT 0.090 268.500 0.700 269.660 ;
        RECT 4.300 268.500 996.660 269.660 ;
        RECT 0.090 262.940 996.660 268.500 ;
        RECT 0.090 261.780 995.700 262.940 ;
        RECT 0.090 259.580 996.660 261.780 ;
        RECT 0.090 258.420 0.700 259.580 ;
        RECT 4.300 258.420 996.660 259.580 ;
        RECT 0.090 252.860 996.660 258.420 ;
        RECT 0.090 251.700 995.700 252.860 ;
        RECT 0.090 249.500 996.660 251.700 ;
        RECT 0.090 248.340 0.700 249.500 ;
        RECT 4.300 248.340 996.660 249.500 ;
        RECT 0.090 242.780 996.660 248.340 ;
        RECT 0.090 241.620 995.700 242.780 ;
        RECT 0.090 239.420 996.660 241.620 ;
        RECT 0.090 238.260 0.700 239.420 ;
        RECT 4.300 238.260 996.660 239.420 ;
        RECT 0.090 232.700 996.660 238.260 ;
        RECT 0.090 231.540 995.700 232.700 ;
        RECT 0.090 229.340 996.660 231.540 ;
        RECT 0.090 228.180 0.700 229.340 ;
        RECT 4.300 228.180 996.660 229.340 ;
        RECT 0.090 222.620 996.660 228.180 ;
        RECT 0.090 221.460 0.700 222.620 ;
        RECT 4.300 221.460 995.700 222.620 ;
        RECT 0.090 212.540 996.660 221.460 ;
        RECT 0.090 211.380 0.700 212.540 ;
        RECT 4.300 211.380 995.700 212.540 ;
        RECT 0.090 205.820 996.660 211.380 ;
        RECT 0.090 204.660 995.700 205.820 ;
        RECT 0.090 202.460 996.660 204.660 ;
        RECT 0.090 201.300 0.700 202.460 ;
        RECT 4.300 201.300 996.660 202.460 ;
        RECT 0.090 195.740 996.660 201.300 ;
        RECT 0.090 194.580 995.700 195.740 ;
        RECT 0.090 192.380 996.660 194.580 ;
        RECT 0.090 191.220 0.700 192.380 ;
        RECT 4.300 191.220 996.660 192.380 ;
        RECT 0.090 185.660 996.660 191.220 ;
        RECT 0.090 184.500 995.700 185.660 ;
        RECT 0.090 182.300 996.660 184.500 ;
        RECT 0.090 181.140 0.700 182.300 ;
        RECT 4.300 181.140 996.660 182.300 ;
        RECT 0.090 175.580 996.660 181.140 ;
        RECT 0.090 174.420 995.700 175.580 ;
        RECT 0.090 172.220 996.660 174.420 ;
        RECT 0.090 171.060 0.700 172.220 ;
        RECT 4.300 171.060 996.660 172.220 ;
        RECT 0.090 165.500 996.660 171.060 ;
        RECT 0.090 164.340 995.700 165.500 ;
        RECT 0.090 162.140 996.660 164.340 ;
        RECT 0.090 160.980 0.700 162.140 ;
        RECT 4.300 160.980 996.660 162.140 ;
        RECT 0.090 155.420 996.660 160.980 ;
        RECT 0.090 154.260 995.700 155.420 ;
        RECT 0.090 152.060 996.660 154.260 ;
        RECT 0.090 150.900 0.700 152.060 ;
        RECT 4.300 150.900 996.660 152.060 ;
        RECT 0.090 145.340 996.660 150.900 ;
        RECT 0.090 144.180 0.700 145.340 ;
        RECT 4.300 144.180 995.700 145.340 ;
        RECT 0.090 135.260 996.660 144.180 ;
        RECT 0.090 134.100 0.700 135.260 ;
        RECT 4.300 134.100 995.700 135.260 ;
        RECT 0.090 128.540 996.660 134.100 ;
        RECT 0.090 127.380 995.700 128.540 ;
        RECT 0.090 125.180 996.660 127.380 ;
        RECT 0.090 124.020 0.700 125.180 ;
        RECT 4.300 124.020 996.660 125.180 ;
        RECT 0.090 118.460 996.660 124.020 ;
        RECT 0.090 117.300 995.700 118.460 ;
        RECT 0.090 115.100 996.660 117.300 ;
        RECT 0.090 113.940 0.700 115.100 ;
        RECT 4.300 113.940 996.660 115.100 ;
        RECT 0.090 108.380 996.660 113.940 ;
        RECT 0.090 107.220 995.700 108.380 ;
        RECT 0.090 105.020 996.660 107.220 ;
        RECT 0.090 103.860 0.700 105.020 ;
        RECT 4.300 103.860 996.660 105.020 ;
        RECT 0.090 98.300 996.660 103.860 ;
        RECT 0.090 97.140 995.700 98.300 ;
        RECT 0.090 94.940 996.660 97.140 ;
        RECT 0.090 93.780 0.700 94.940 ;
        RECT 4.300 93.780 996.660 94.940 ;
        RECT 0.090 88.220 996.660 93.780 ;
        RECT 0.090 87.060 995.700 88.220 ;
        RECT 0.090 84.860 996.660 87.060 ;
        RECT 0.090 83.700 0.700 84.860 ;
        RECT 4.300 83.700 996.660 84.860 ;
        RECT 0.090 78.140 996.660 83.700 ;
        RECT 0.090 76.980 995.700 78.140 ;
        RECT 0.090 74.780 996.660 76.980 ;
        RECT 0.090 73.620 0.700 74.780 ;
        RECT 4.300 73.620 996.660 74.780 ;
        RECT 0.090 68.060 996.660 73.620 ;
        RECT 0.090 66.900 0.700 68.060 ;
        RECT 4.300 66.900 995.700 68.060 ;
        RECT 0.090 57.980 996.660 66.900 ;
        RECT 0.090 56.820 0.700 57.980 ;
        RECT 4.300 56.820 995.700 57.980 ;
        RECT 0.090 51.260 996.660 56.820 ;
        RECT 0.090 50.100 995.700 51.260 ;
        RECT 0.090 47.900 996.660 50.100 ;
        RECT 0.090 46.740 0.700 47.900 ;
        RECT 4.300 46.740 996.660 47.900 ;
        RECT 0.090 41.180 996.660 46.740 ;
        RECT 0.090 40.020 995.700 41.180 ;
        RECT 0.090 37.820 996.660 40.020 ;
        RECT 0.090 36.660 0.700 37.820 ;
        RECT 4.300 36.660 996.660 37.820 ;
        RECT 0.090 31.100 996.660 36.660 ;
        RECT 0.090 29.940 995.700 31.100 ;
        RECT 0.090 27.740 996.660 29.940 ;
        RECT 0.090 26.580 0.700 27.740 ;
        RECT 4.300 26.580 996.660 27.740 ;
        RECT 0.090 21.020 996.660 26.580 ;
        RECT 0.090 19.860 995.700 21.020 ;
        RECT 0.090 17.660 996.660 19.860 ;
        RECT 0.090 16.500 0.700 17.660 ;
        RECT 4.300 16.500 996.660 17.660 ;
        RECT 0.090 10.940 996.660 16.500 ;
        RECT 0.090 9.780 995.700 10.940 ;
        RECT 0.090 7.580 996.660 9.780 ;
        RECT 0.090 6.860 0.700 7.580 ;
        RECT 4.300 6.860 996.660 7.580 ;
      LAYER Metal4 ;
        RECT 11.900 17.450 21.940 982.710 ;
        RECT 24.140 17.450 98.740 982.710 ;
        RECT 100.940 17.450 175.540 982.710 ;
        RECT 177.740 17.450 252.340 982.710 ;
        RECT 254.540 17.450 329.140 982.710 ;
        RECT 331.340 17.450 405.940 982.710 ;
        RECT 408.140 17.450 482.740 982.710 ;
        RECT 484.940 17.450 559.540 982.710 ;
        RECT 561.740 17.450 636.340 982.710 ;
        RECT 638.540 17.450 713.140 982.710 ;
        RECT 715.340 17.450 789.940 982.710 ;
        RECT 792.140 17.450 866.740 982.710 ;
        RECT 868.940 17.450 870.660 982.710 ;
      LAYER Metal5 ;
        RECT 11.820 75.660 799.060 696.020 ;
  END
END caravel_hack_soc
END LIBRARY

