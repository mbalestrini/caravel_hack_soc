magic
tech gf180mcuC
magscale 1 5
timestamp 1670275738
<< obsm1 >>
rect 672 855 59304 58729
<< metal2 >>
rect 0 59600 56 59900
rect 672 59600 728 59900
rect 1008 59600 1064 59900
rect 1680 59600 1736 59900
rect 2352 59600 2408 59900
rect 3024 59600 3080 59900
rect 3360 59600 3416 59900
rect 4032 59600 4088 59900
rect 4704 59600 4760 59900
rect 5040 59600 5096 59900
rect 5712 59600 5768 59900
rect 6384 59600 6440 59900
rect 7056 59600 7112 59900
rect 7392 59600 7448 59900
rect 8064 59600 8120 59900
rect 8736 59600 8792 59900
rect 9408 59600 9464 59900
rect 9744 59600 9800 59900
rect 10416 59600 10472 59900
rect 11088 59600 11144 59900
rect 11424 59600 11480 59900
rect 12096 59600 12152 59900
rect 12768 59600 12824 59900
rect 13440 59600 13496 59900
rect 13776 59600 13832 59900
rect 14448 59600 14504 59900
rect 15120 59600 15176 59900
rect 15792 59600 15848 59900
rect 16128 59600 16184 59900
rect 16800 59600 16856 59900
rect 17472 59600 17528 59900
rect 17808 59600 17864 59900
rect 18480 59600 18536 59900
rect 19152 59600 19208 59900
rect 19824 59600 19880 59900
rect 20160 59600 20216 59900
rect 20832 59600 20888 59900
rect 21504 59600 21560 59900
rect 21840 59600 21896 59900
rect 22512 59600 22568 59900
rect 23184 59600 23240 59900
rect 23856 59600 23912 59900
rect 24192 59600 24248 59900
rect 24864 59600 24920 59900
rect 25536 59600 25592 59900
rect 26208 59600 26264 59900
rect 26544 59600 26600 59900
rect 27216 59600 27272 59900
rect 27888 59600 27944 59900
rect 28224 59600 28280 59900
rect 28896 59600 28952 59900
rect 29568 59600 29624 59900
rect 30240 59600 30296 59900
rect 30576 59600 30632 59900
rect 31248 59600 31304 59900
rect 31920 59600 31976 59900
rect 32592 59600 32648 59900
rect 32928 59600 32984 59900
rect 33600 59600 33656 59900
rect 34272 59600 34328 59900
rect 34608 59600 34664 59900
rect 35280 59600 35336 59900
rect 35952 59600 36008 59900
rect 36624 59600 36680 59900
rect 36960 59600 37016 59900
rect 37632 59600 37688 59900
rect 38304 59600 38360 59900
rect 38976 59600 39032 59900
rect 39312 59600 39368 59900
rect 39984 59600 40040 59900
rect 40656 59600 40712 59900
rect 40992 59600 41048 59900
rect 41664 59600 41720 59900
rect 42336 59600 42392 59900
rect 43008 59600 43064 59900
rect 43344 59600 43400 59900
rect 44016 59600 44072 59900
rect 44688 59600 44744 59900
rect 45360 59600 45416 59900
rect 45696 59600 45752 59900
rect 46368 59600 46424 59900
rect 47040 59600 47096 59900
rect 47376 59600 47432 59900
rect 48048 59600 48104 59900
rect 48720 59600 48776 59900
rect 49392 59600 49448 59900
rect 49728 59600 49784 59900
rect 50400 59600 50456 59900
rect 51072 59600 51128 59900
rect 51408 59600 51464 59900
rect 52080 59600 52136 59900
rect 52752 59600 52808 59900
rect 53424 59600 53480 59900
rect 53760 59600 53816 59900
rect 54432 59600 54488 59900
rect 55104 59600 55160 59900
rect 55776 59600 55832 59900
rect 56112 59600 56168 59900
rect 56784 59600 56840 59900
rect 57456 59600 57512 59900
rect 57792 59600 57848 59900
rect 58464 59600 58520 59900
rect 59136 59600 59192 59900
rect 59808 59600 59864 59900
rect 0 100 56 400
rect 336 100 392 400
rect 1008 100 1064 400
rect 1680 100 1736 400
rect 2016 100 2072 400
rect 2688 100 2744 400
rect 3360 100 3416 400
rect 4032 100 4088 400
rect 4368 100 4424 400
rect 5040 100 5096 400
rect 5712 100 5768 400
rect 6048 100 6104 400
rect 6720 100 6776 400
rect 7392 100 7448 400
rect 8064 100 8120 400
rect 8400 100 8456 400
rect 9072 100 9128 400
rect 9744 100 9800 400
rect 10416 100 10472 400
rect 10752 100 10808 400
rect 11424 100 11480 400
rect 12096 100 12152 400
rect 12432 100 12488 400
rect 13104 100 13160 400
rect 13776 100 13832 400
rect 14448 100 14504 400
rect 14784 100 14840 400
rect 15456 100 15512 400
rect 16128 100 16184 400
rect 16800 100 16856 400
rect 17136 100 17192 400
rect 17808 100 17864 400
rect 18480 100 18536 400
rect 18816 100 18872 400
rect 19488 100 19544 400
rect 20160 100 20216 400
rect 20832 100 20888 400
rect 21168 100 21224 400
rect 21840 100 21896 400
rect 22512 100 22568 400
rect 23184 100 23240 400
rect 23520 100 23576 400
rect 24192 100 24248 400
rect 24864 100 24920 400
rect 25200 100 25256 400
rect 25872 100 25928 400
rect 26544 100 26600 400
rect 27216 100 27272 400
rect 27552 100 27608 400
rect 28224 100 28280 400
rect 28896 100 28952 400
rect 29232 100 29288 400
rect 29904 100 29960 400
rect 30576 100 30632 400
rect 31248 100 31304 400
rect 31584 100 31640 400
rect 32256 100 32312 400
rect 32928 100 32984 400
rect 33600 100 33656 400
rect 33936 100 33992 400
rect 34608 100 34664 400
rect 35280 100 35336 400
rect 35616 100 35672 400
rect 36288 100 36344 400
rect 36960 100 37016 400
rect 37632 100 37688 400
rect 37968 100 38024 400
rect 38640 100 38696 400
rect 39312 100 39368 400
rect 39984 100 40040 400
rect 40320 100 40376 400
rect 40992 100 41048 400
rect 41664 100 41720 400
rect 42000 100 42056 400
rect 42672 100 42728 400
rect 43344 100 43400 400
rect 44016 100 44072 400
rect 44352 100 44408 400
rect 45024 100 45080 400
rect 45696 100 45752 400
rect 46368 100 46424 400
rect 46704 100 46760 400
rect 47376 100 47432 400
rect 48048 100 48104 400
rect 48384 100 48440 400
rect 49056 100 49112 400
rect 49728 100 49784 400
rect 50400 100 50456 400
rect 50736 100 50792 400
rect 51408 100 51464 400
rect 52080 100 52136 400
rect 52752 100 52808 400
rect 53088 100 53144 400
rect 53760 100 53816 400
rect 54432 100 54488 400
rect 54768 100 54824 400
rect 55440 100 55496 400
rect 56112 100 56168 400
rect 56784 100 56840 400
rect 57120 100 57176 400
rect 57792 100 57848 400
rect 58464 100 58520 400
rect 58800 100 58856 400
rect 59472 100 59528 400
<< obsm2 >>
rect 86 59570 642 59631
rect 758 59570 978 59631
rect 1094 59570 1650 59631
rect 1766 59570 2322 59631
rect 2438 59570 2994 59631
rect 3110 59570 3330 59631
rect 3446 59570 4002 59631
rect 4118 59570 4674 59631
rect 4790 59570 5010 59631
rect 5126 59570 5682 59631
rect 5798 59570 6354 59631
rect 6470 59570 7026 59631
rect 7142 59570 7362 59631
rect 7478 59570 8034 59631
rect 8150 59570 8706 59631
rect 8822 59570 9378 59631
rect 9494 59570 9714 59631
rect 9830 59570 10386 59631
rect 10502 59570 11058 59631
rect 11174 59570 11394 59631
rect 11510 59570 12066 59631
rect 12182 59570 12738 59631
rect 12854 59570 13410 59631
rect 13526 59570 13746 59631
rect 13862 59570 14418 59631
rect 14534 59570 15090 59631
rect 15206 59570 15762 59631
rect 15878 59570 16098 59631
rect 16214 59570 16770 59631
rect 16886 59570 17442 59631
rect 17558 59570 17778 59631
rect 17894 59570 18450 59631
rect 18566 59570 19122 59631
rect 19238 59570 19794 59631
rect 19910 59570 20130 59631
rect 20246 59570 20802 59631
rect 20918 59570 21474 59631
rect 21590 59570 21810 59631
rect 21926 59570 22482 59631
rect 22598 59570 23154 59631
rect 23270 59570 23826 59631
rect 23942 59570 24162 59631
rect 24278 59570 24834 59631
rect 24950 59570 25506 59631
rect 25622 59570 26178 59631
rect 26294 59570 26514 59631
rect 26630 59570 27186 59631
rect 27302 59570 27858 59631
rect 27974 59570 28194 59631
rect 28310 59570 28866 59631
rect 28982 59570 29538 59631
rect 29654 59570 30210 59631
rect 30326 59570 30546 59631
rect 30662 59570 31218 59631
rect 31334 59570 31890 59631
rect 32006 59570 32562 59631
rect 32678 59570 32898 59631
rect 33014 59570 33570 59631
rect 33686 59570 34242 59631
rect 34358 59570 34578 59631
rect 34694 59570 35250 59631
rect 35366 59570 35922 59631
rect 36038 59570 36594 59631
rect 36710 59570 36930 59631
rect 37046 59570 37602 59631
rect 37718 59570 38274 59631
rect 38390 59570 38946 59631
rect 39062 59570 39282 59631
rect 39398 59570 39954 59631
rect 40070 59570 40626 59631
rect 40742 59570 40962 59631
rect 41078 59570 41634 59631
rect 41750 59570 42306 59631
rect 42422 59570 42978 59631
rect 43094 59570 43314 59631
rect 43430 59570 43986 59631
rect 44102 59570 44658 59631
rect 44774 59570 45330 59631
rect 45446 59570 45666 59631
rect 45782 59570 46338 59631
rect 46454 59570 47010 59631
rect 47126 59570 47346 59631
rect 47462 59570 48018 59631
rect 48134 59570 48690 59631
rect 48806 59570 49362 59631
rect 49478 59570 49698 59631
rect 49814 59570 50370 59631
rect 50486 59570 51042 59631
rect 51158 59570 51378 59631
rect 51494 59570 52050 59631
rect 52166 59570 52722 59631
rect 52838 59570 53394 59631
rect 53510 59570 53730 59631
rect 53846 59570 54402 59631
rect 54518 59570 55074 59631
rect 55190 59570 55746 59631
rect 55862 59570 56082 59631
rect 56198 59570 56754 59631
rect 56870 59570 57426 59631
rect 57542 59570 57762 59631
rect 57878 59570 58434 59631
rect 58550 59570 59106 59631
rect 14 430 59178 59570
rect 86 400 306 430
rect 422 400 978 430
rect 1094 400 1650 430
rect 1766 400 1986 430
rect 2102 400 2658 430
rect 2774 400 3330 430
rect 3446 400 4002 430
rect 4118 400 4338 430
rect 4454 400 5010 430
rect 5126 400 5682 430
rect 5798 400 6018 430
rect 6134 400 6690 430
rect 6806 400 7362 430
rect 7478 400 8034 430
rect 8150 400 8370 430
rect 8486 400 9042 430
rect 9158 400 9714 430
rect 9830 400 10386 430
rect 10502 400 10722 430
rect 10838 400 11394 430
rect 11510 400 12066 430
rect 12182 400 12402 430
rect 12518 400 13074 430
rect 13190 400 13746 430
rect 13862 400 14418 430
rect 14534 400 14754 430
rect 14870 400 15426 430
rect 15542 400 16098 430
rect 16214 400 16770 430
rect 16886 400 17106 430
rect 17222 400 17778 430
rect 17894 400 18450 430
rect 18566 400 18786 430
rect 18902 400 19458 430
rect 19574 400 20130 430
rect 20246 400 20802 430
rect 20918 400 21138 430
rect 21254 400 21810 430
rect 21926 400 22482 430
rect 22598 400 23154 430
rect 23270 400 23490 430
rect 23606 400 24162 430
rect 24278 400 24834 430
rect 24950 400 25170 430
rect 25286 400 25842 430
rect 25958 400 26514 430
rect 26630 400 27186 430
rect 27302 400 27522 430
rect 27638 400 28194 430
rect 28310 400 28866 430
rect 28982 400 29202 430
rect 29318 400 29874 430
rect 29990 400 30546 430
rect 30662 400 31218 430
rect 31334 400 31554 430
rect 31670 400 32226 430
rect 32342 400 32898 430
rect 33014 400 33570 430
rect 33686 400 33906 430
rect 34022 400 34578 430
rect 34694 400 35250 430
rect 35366 400 35586 430
rect 35702 400 36258 430
rect 36374 400 36930 430
rect 37046 400 37602 430
rect 37718 400 37938 430
rect 38054 400 38610 430
rect 38726 400 39282 430
rect 39398 400 39954 430
rect 40070 400 40290 430
rect 40406 400 40962 430
rect 41078 400 41634 430
rect 41750 400 41970 430
rect 42086 400 42642 430
rect 42758 400 43314 430
rect 43430 400 43986 430
rect 44102 400 44322 430
rect 44438 400 44994 430
rect 45110 400 45666 430
rect 45782 400 46338 430
rect 46454 400 46674 430
rect 46790 400 47346 430
rect 47462 400 48018 430
rect 48134 400 48354 430
rect 48470 400 49026 430
rect 49142 400 49698 430
rect 49814 400 50370 430
rect 50486 400 50706 430
rect 50822 400 51378 430
rect 51494 400 52050 430
rect 52166 400 52722 430
rect 52838 400 53058 430
rect 53174 400 53730 430
rect 53846 400 54402 430
rect 54518 400 54738 430
rect 54854 400 55410 430
rect 55526 400 56082 430
rect 56198 400 56754 430
rect 56870 400 57090 430
rect 57206 400 57762 430
rect 57878 400 58434 430
rect 58550 400 58770 430
rect 58886 400 59178 430
<< metal3 >>
rect 59600 59808 59900 59864
rect 100 59472 400 59528
rect 59600 59136 59900 59192
rect 100 58800 400 58856
rect 100 58464 400 58520
rect 59600 58464 59900 58520
rect 100 57792 400 57848
rect 59600 57792 59900 57848
rect 59600 57456 59900 57512
rect 100 57120 400 57176
rect 100 56784 400 56840
rect 59600 56784 59900 56840
rect 100 56112 400 56168
rect 59600 56112 59900 56168
rect 59600 55776 59900 55832
rect 100 55440 400 55496
rect 59600 55104 59900 55160
rect 100 54768 400 54824
rect 100 54432 400 54488
rect 59600 54432 59900 54488
rect 100 53760 400 53816
rect 59600 53760 59900 53816
rect 59600 53424 59900 53480
rect 100 53088 400 53144
rect 100 52752 400 52808
rect 59600 52752 59900 52808
rect 100 52080 400 52136
rect 59600 52080 59900 52136
rect 100 51408 400 51464
rect 59600 51408 59900 51464
rect 59600 51072 59900 51128
rect 100 50736 400 50792
rect 100 50400 400 50456
rect 59600 50400 59900 50456
rect 100 49728 400 49784
rect 59600 49728 59900 49784
rect 59600 49392 59900 49448
rect 100 49056 400 49112
rect 59600 48720 59900 48776
rect 100 48384 400 48440
rect 100 48048 400 48104
rect 59600 48048 59900 48104
rect 100 47376 400 47432
rect 59600 47376 59900 47432
rect 59600 47040 59900 47096
rect 100 46704 400 46760
rect 100 46368 400 46424
rect 59600 46368 59900 46424
rect 100 45696 400 45752
rect 59600 45696 59900 45752
rect 59600 45360 59900 45416
rect 100 45024 400 45080
rect 59600 44688 59900 44744
rect 100 44352 400 44408
rect 100 44016 400 44072
rect 59600 44016 59900 44072
rect 100 43344 400 43400
rect 59600 43344 59900 43400
rect 59600 43008 59900 43064
rect 100 42672 400 42728
rect 59600 42336 59900 42392
rect 100 42000 400 42056
rect 100 41664 400 41720
rect 59600 41664 59900 41720
rect 100 40992 400 41048
rect 59600 40992 59900 41048
rect 59600 40656 59900 40712
rect 100 40320 400 40376
rect 100 39984 400 40040
rect 59600 39984 59900 40040
rect 100 39312 400 39368
rect 59600 39312 59900 39368
rect 59600 38976 59900 39032
rect 100 38640 400 38696
rect 59600 38304 59900 38360
rect 100 37968 400 38024
rect 100 37632 400 37688
rect 59600 37632 59900 37688
rect 100 36960 400 37016
rect 59600 36960 59900 37016
rect 59600 36624 59900 36680
rect 100 36288 400 36344
rect 59600 35952 59900 36008
rect 100 35616 400 35672
rect 100 35280 400 35336
rect 59600 35280 59900 35336
rect 100 34608 400 34664
rect 59600 34608 59900 34664
rect 59600 34272 59900 34328
rect 100 33936 400 33992
rect 100 33600 400 33656
rect 59600 33600 59900 33656
rect 100 32928 400 32984
rect 59600 32928 59900 32984
rect 59600 32592 59900 32648
rect 100 32256 400 32312
rect 59600 31920 59900 31976
rect 100 31584 400 31640
rect 100 31248 400 31304
rect 59600 31248 59900 31304
rect 100 30576 400 30632
rect 59600 30576 59900 30632
rect 59600 30240 59900 30296
rect 100 29904 400 29960
rect 59600 29568 59900 29624
rect 100 29232 400 29288
rect 100 28896 400 28952
rect 59600 28896 59900 28952
rect 100 28224 400 28280
rect 59600 28224 59900 28280
rect 59600 27888 59900 27944
rect 100 27552 400 27608
rect 100 27216 400 27272
rect 59600 27216 59900 27272
rect 100 26544 400 26600
rect 59600 26544 59900 26600
rect 59600 26208 59900 26264
rect 100 25872 400 25928
rect 59600 25536 59900 25592
rect 100 25200 400 25256
rect 100 24864 400 24920
rect 59600 24864 59900 24920
rect 100 24192 400 24248
rect 59600 24192 59900 24248
rect 59600 23856 59900 23912
rect 100 23520 400 23576
rect 100 23184 400 23240
rect 59600 23184 59900 23240
rect 100 22512 400 22568
rect 59600 22512 59900 22568
rect 100 21840 400 21896
rect 59600 21840 59900 21896
rect 59600 21504 59900 21560
rect 100 21168 400 21224
rect 100 20832 400 20888
rect 59600 20832 59900 20888
rect 100 20160 400 20216
rect 59600 20160 59900 20216
rect 59600 19824 59900 19880
rect 100 19488 400 19544
rect 59600 19152 59900 19208
rect 100 18816 400 18872
rect 100 18480 400 18536
rect 59600 18480 59900 18536
rect 100 17808 400 17864
rect 59600 17808 59900 17864
rect 59600 17472 59900 17528
rect 100 17136 400 17192
rect 100 16800 400 16856
rect 59600 16800 59900 16856
rect 100 16128 400 16184
rect 59600 16128 59900 16184
rect 59600 15792 59900 15848
rect 100 15456 400 15512
rect 59600 15120 59900 15176
rect 100 14784 400 14840
rect 100 14448 400 14504
rect 59600 14448 59900 14504
rect 100 13776 400 13832
rect 59600 13776 59900 13832
rect 59600 13440 59900 13496
rect 100 13104 400 13160
rect 59600 12768 59900 12824
rect 100 12432 400 12488
rect 100 12096 400 12152
rect 59600 12096 59900 12152
rect 100 11424 400 11480
rect 59600 11424 59900 11480
rect 59600 11088 59900 11144
rect 100 10752 400 10808
rect 100 10416 400 10472
rect 59600 10416 59900 10472
rect 100 9744 400 9800
rect 59600 9744 59900 9800
rect 59600 9408 59900 9464
rect 100 9072 400 9128
rect 59600 8736 59900 8792
rect 100 8400 400 8456
rect 100 8064 400 8120
rect 59600 8064 59900 8120
rect 100 7392 400 7448
rect 59600 7392 59900 7448
rect 59600 7056 59900 7112
rect 100 6720 400 6776
rect 59600 6384 59900 6440
rect 100 6048 400 6104
rect 100 5712 400 5768
rect 59600 5712 59900 5768
rect 100 5040 400 5096
rect 59600 5040 59900 5096
rect 59600 4704 59900 4760
rect 100 4368 400 4424
rect 100 4032 400 4088
rect 59600 4032 59900 4088
rect 100 3360 400 3416
rect 59600 3360 59900 3416
rect 59600 3024 59900 3080
rect 100 2688 400 2744
rect 59600 2352 59900 2408
rect 100 2016 400 2072
rect 100 1680 400 1736
rect 59600 1680 59900 1736
rect 100 1008 400 1064
rect 59600 1008 59900 1064
rect 59600 672 59900 728
rect 100 336 400 392
rect 59600 0 59900 56
<< obsm3 >>
rect 9 59778 59570 59850
rect 9 59558 59682 59778
rect 9 59442 70 59558
rect 430 59442 59682 59558
rect 9 59222 59682 59442
rect 9 59106 59570 59222
rect 9 58886 59682 59106
rect 9 58770 70 58886
rect 430 58770 59682 58886
rect 9 58550 59682 58770
rect 9 58434 70 58550
rect 430 58434 59570 58550
rect 9 57878 59682 58434
rect 9 57762 70 57878
rect 430 57762 59570 57878
rect 9 57542 59682 57762
rect 9 57426 59570 57542
rect 9 57206 59682 57426
rect 9 57090 70 57206
rect 430 57090 59682 57206
rect 9 56870 59682 57090
rect 9 56754 70 56870
rect 430 56754 59570 56870
rect 9 56198 59682 56754
rect 9 56082 70 56198
rect 430 56082 59570 56198
rect 9 55862 59682 56082
rect 9 55746 59570 55862
rect 9 55526 59682 55746
rect 9 55410 70 55526
rect 430 55410 59682 55526
rect 9 55190 59682 55410
rect 9 55074 59570 55190
rect 9 54854 59682 55074
rect 9 54738 70 54854
rect 430 54738 59682 54854
rect 9 54518 59682 54738
rect 9 54402 70 54518
rect 430 54402 59570 54518
rect 9 53846 59682 54402
rect 9 53730 70 53846
rect 430 53730 59570 53846
rect 9 53510 59682 53730
rect 9 53394 59570 53510
rect 9 53174 59682 53394
rect 9 53058 70 53174
rect 430 53058 59682 53174
rect 9 52838 59682 53058
rect 9 52722 70 52838
rect 430 52722 59570 52838
rect 9 52166 59682 52722
rect 9 52050 70 52166
rect 430 52050 59570 52166
rect 9 51494 59682 52050
rect 9 51378 70 51494
rect 430 51378 59570 51494
rect 9 51158 59682 51378
rect 9 51042 59570 51158
rect 9 50822 59682 51042
rect 9 50706 70 50822
rect 430 50706 59682 50822
rect 9 50486 59682 50706
rect 9 50370 70 50486
rect 430 50370 59570 50486
rect 9 49814 59682 50370
rect 9 49698 70 49814
rect 430 49698 59570 49814
rect 9 49478 59682 49698
rect 9 49362 59570 49478
rect 9 49142 59682 49362
rect 9 49026 70 49142
rect 430 49026 59682 49142
rect 9 48806 59682 49026
rect 9 48690 59570 48806
rect 9 48470 59682 48690
rect 9 48354 70 48470
rect 430 48354 59682 48470
rect 9 48134 59682 48354
rect 9 48018 70 48134
rect 430 48018 59570 48134
rect 9 47462 59682 48018
rect 9 47346 70 47462
rect 430 47346 59570 47462
rect 9 47126 59682 47346
rect 9 47010 59570 47126
rect 9 46790 59682 47010
rect 9 46674 70 46790
rect 430 46674 59682 46790
rect 9 46454 59682 46674
rect 9 46338 70 46454
rect 430 46338 59570 46454
rect 9 45782 59682 46338
rect 9 45666 70 45782
rect 430 45666 59570 45782
rect 9 45446 59682 45666
rect 9 45330 59570 45446
rect 9 45110 59682 45330
rect 9 44994 70 45110
rect 430 44994 59682 45110
rect 9 44774 59682 44994
rect 9 44658 59570 44774
rect 9 44438 59682 44658
rect 9 44322 70 44438
rect 430 44322 59682 44438
rect 9 44102 59682 44322
rect 9 43986 70 44102
rect 430 43986 59570 44102
rect 9 43430 59682 43986
rect 9 43314 70 43430
rect 430 43314 59570 43430
rect 9 43094 59682 43314
rect 9 42978 59570 43094
rect 9 42758 59682 42978
rect 9 42642 70 42758
rect 430 42642 59682 42758
rect 9 42422 59682 42642
rect 9 42306 59570 42422
rect 9 42086 59682 42306
rect 9 41970 70 42086
rect 430 41970 59682 42086
rect 9 41750 59682 41970
rect 9 41634 70 41750
rect 430 41634 59570 41750
rect 9 41078 59682 41634
rect 9 40962 70 41078
rect 430 40962 59570 41078
rect 9 40742 59682 40962
rect 9 40626 59570 40742
rect 9 40406 59682 40626
rect 9 40290 70 40406
rect 430 40290 59682 40406
rect 9 40070 59682 40290
rect 9 39954 70 40070
rect 430 39954 59570 40070
rect 9 39398 59682 39954
rect 9 39282 70 39398
rect 430 39282 59570 39398
rect 9 39062 59682 39282
rect 9 38946 59570 39062
rect 9 38726 59682 38946
rect 9 38610 70 38726
rect 430 38610 59682 38726
rect 9 38390 59682 38610
rect 9 38274 59570 38390
rect 9 38054 59682 38274
rect 9 37938 70 38054
rect 430 37938 59682 38054
rect 9 37718 59682 37938
rect 9 37602 70 37718
rect 430 37602 59570 37718
rect 9 37046 59682 37602
rect 9 36930 70 37046
rect 430 36930 59570 37046
rect 9 36710 59682 36930
rect 9 36594 59570 36710
rect 9 36374 59682 36594
rect 9 36258 70 36374
rect 430 36258 59682 36374
rect 9 36038 59682 36258
rect 9 35922 59570 36038
rect 9 35702 59682 35922
rect 9 35586 70 35702
rect 430 35586 59682 35702
rect 9 35366 59682 35586
rect 9 35250 70 35366
rect 430 35250 59570 35366
rect 9 34694 59682 35250
rect 9 34578 70 34694
rect 430 34578 59570 34694
rect 9 34358 59682 34578
rect 9 34242 59570 34358
rect 9 34022 59682 34242
rect 9 33906 70 34022
rect 430 33906 59682 34022
rect 9 33686 59682 33906
rect 9 33570 70 33686
rect 430 33570 59570 33686
rect 9 33014 59682 33570
rect 9 32898 70 33014
rect 430 32898 59570 33014
rect 9 32678 59682 32898
rect 9 32562 59570 32678
rect 9 32342 59682 32562
rect 9 32226 70 32342
rect 430 32226 59682 32342
rect 9 32006 59682 32226
rect 9 31890 59570 32006
rect 9 31670 59682 31890
rect 9 31554 70 31670
rect 430 31554 59682 31670
rect 9 31334 59682 31554
rect 9 31218 70 31334
rect 430 31218 59570 31334
rect 9 30662 59682 31218
rect 9 30546 70 30662
rect 430 30546 59570 30662
rect 9 30326 59682 30546
rect 9 30210 59570 30326
rect 9 29990 59682 30210
rect 9 29874 70 29990
rect 430 29874 59682 29990
rect 9 29654 59682 29874
rect 9 29538 59570 29654
rect 9 29318 59682 29538
rect 9 29202 70 29318
rect 430 29202 59682 29318
rect 9 28982 59682 29202
rect 9 28866 70 28982
rect 430 28866 59570 28982
rect 9 28310 59682 28866
rect 9 28194 70 28310
rect 430 28194 59570 28310
rect 9 27974 59682 28194
rect 9 27858 59570 27974
rect 9 27638 59682 27858
rect 9 27522 70 27638
rect 430 27522 59682 27638
rect 9 27302 59682 27522
rect 9 27186 70 27302
rect 430 27186 59570 27302
rect 9 26630 59682 27186
rect 9 26514 70 26630
rect 430 26514 59570 26630
rect 9 26294 59682 26514
rect 9 26178 59570 26294
rect 9 25958 59682 26178
rect 9 25842 70 25958
rect 430 25842 59682 25958
rect 9 25622 59682 25842
rect 9 25506 59570 25622
rect 9 25286 59682 25506
rect 9 25170 70 25286
rect 430 25170 59682 25286
rect 9 24950 59682 25170
rect 9 24834 70 24950
rect 430 24834 59570 24950
rect 9 24278 59682 24834
rect 9 24162 70 24278
rect 430 24162 59570 24278
rect 9 23942 59682 24162
rect 9 23826 59570 23942
rect 9 23606 59682 23826
rect 9 23490 70 23606
rect 430 23490 59682 23606
rect 9 23270 59682 23490
rect 9 23154 70 23270
rect 430 23154 59570 23270
rect 9 22598 59682 23154
rect 9 22482 70 22598
rect 430 22482 59570 22598
rect 9 21926 59682 22482
rect 9 21810 70 21926
rect 430 21810 59570 21926
rect 9 21590 59682 21810
rect 9 21474 59570 21590
rect 9 21254 59682 21474
rect 9 21138 70 21254
rect 430 21138 59682 21254
rect 9 20918 59682 21138
rect 9 20802 70 20918
rect 430 20802 59570 20918
rect 9 20246 59682 20802
rect 9 20130 70 20246
rect 430 20130 59570 20246
rect 9 19910 59682 20130
rect 9 19794 59570 19910
rect 9 19574 59682 19794
rect 9 19458 70 19574
rect 430 19458 59682 19574
rect 9 19238 59682 19458
rect 9 19122 59570 19238
rect 9 18902 59682 19122
rect 9 18786 70 18902
rect 430 18786 59682 18902
rect 9 18566 59682 18786
rect 9 18450 70 18566
rect 430 18450 59570 18566
rect 9 17894 59682 18450
rect 9 17778 70 17894
rect 430 17778 59570 17894
rect 9 17558 59682 17778
rect 9 17442 59570 17558
rect 9 17222 59682 17442
rect 9 17106 70 17222
rect 430 17106 59682 17222
rect 9 16886 59682 17106
rect 9 16770 70 16886
rect 430 16770 59570 16886
rect 9 16214 59682 16770
rect 9 16098 70 16214
rect 430 16098 59570 16214
rect 9 15878 59682 16098
rect 9 15762 59570 15878
rect 9 15542 59682 15762
rect 9 15426 70 15542
rect 430 15426 59682 15542
rect 9 15206 59682 15426
rect 9 15090 59570 15206
rect 9 14870 59682 15090
rect 9 14754 70 14870
rect 430 14754 59682 14870
rect 9 14534 59682 14754
rect 9 14418 70 14534
rect 430 14418 59570 14534
rect 9 13862 59682 14418
rect 9 13746 70 13862
rect 430 13746 59570 13862
rect 9 13526 59682 13746
rect 9 13410 59570 13526
rect 9 13190 59682 13410
rect 9 13074 70 13190
rect 430 13074 59682 13190
rect 9 12854 59682 13074
rect 9 12738 59570 12854
rect 9 12518 59682 12738
rect 9 12402 70 12518
rect 430 12402 59682 12518
rect 9 12182 59682 12402
rect 9 12066 70 12182
rect 430 12066 59570 12182
rect 9 11510 59682 12066
rect 9 11394 70 11510
rect 430 11394 59570 11510
rect 9 11174 59682 11394
rect 9 11058 59570 11174
rect 9 10838 59682 11058
rect 9 10722 70 10838
rect 430 10722 59682 10838
rect 9 10502 59682 10722
rect 9 10386 70 10502
rect 430 10386 59570 10502
rect 9 9830 59682 10386
rect 9 9714 70 9830
rect 430 9714 59570 9830
rect 9 9494 59682 9714
rect 9 9378 59570 9494
rect 9 9158 59682 9378
rect 9 9042 70 9158
rect 430 9042 59682 9158
rect 9 8822 59682 9042
rect 9 8706 59570 8822
rect 9 8486 59682 8706
rect 9 8370 70 8486
rect 430 8370 59682 8486
rect 9 8150 59682 8370
rect 9 8034 70 8150
rect 430 8034 59570 8150
rect 9 7478 59682 8034
rect 9 7362 70 7478
rect 430 7362 59570 7478
rect 9 7142 59682 7362
rect 9 7026 59570 7142
rect 9 6806 59682 7026
rect 9 6690 70 6806
rect 430 6690 59682 6806
rect 9 6470 59682 6690
rect 9 6354 59570 6470
rect 9 6134 59682 6354
rect 9 6018 70 6134
rect 430 6018 59682 6134
rect 9 5798 59682 6018
rect 9 5682 70 5798
rect 430 5682 59570 5798
rect 9 5126 59682 5682
rect 9 5010 70 5126
rect 430 5010 59570 5126
rect 9 4790 59682 5010
rect 9 4674 59570 4790
rect 9 4454 59682 4674
rect 9 4338 70 4454
rect 430 4338 59682 4454
rect 9 4118 59682 4338
rect 9 4002 70 4118
rect 430 4002 59570 4118
rect 9 3446 59682 4002
rect 9 3330 70 3446
rect 430 3330 59570 3446
rect 9 3110 59682 3330
rect 9 2994 59570 3110
rect 9 2774 59682 2994
rect 9 2658 70 2774
rect 430 2658 59682 2774
rect 9 2438 59682 2658
rect 9 2322 59570 2438
rect 9 2102 59682 2322
rect 9 1986 70 2102
rect 430 1986 59682 2102
rect 9 1766 59682 1986
rect 9 1650 70 1766
rect 430 1650 59570 1766
rect 9 1094 59682 1650
rect 9 978 70 1094
rect 430 978 59570 1094
rect 9 758 59682 978
rect 9 642 59570 758
rect 9 422 59682 642
rect 9 350 70 422
rect 430 350 59682 422
<< metal4 >>
rect 2224 1538 2384 58438
rect 9904 1538 10064 58438
rect 17584 1538 17744 58438
rect 25264 1538 25424 58438
rect 32944 1538 33104 58438
rect 40624 1538 40784 58438
rect 48304 1538 48464 58438
rect 55984 1538 56144 58438
<< obsm4 >>
rect 1246 1745 2194 58231
rect 2414 1745 9874 58231
rect 10094 1745 17554 58231
rect 17774 1745 25234 58231
rect 25454 1745 32914 58231
rect 33134 1745 40594 58231
rect 40814 1745 48274 58231
rect 48494 1745 54922 58231
<< obsm5 >>
rect 1238 9862 47706 48826
<< labels >>
rlabel metal3 s 100 20832 400 20888 6 io_in[0]
port 1 nsew signal input
rlabel metal3 s 100 27552 400 27608 6 io_in[10]
port 2 nsew signal input
rlabel metal3 s 100 24864 400 24920 6 io_in[11]
port 3 nsew signal input
rlabel metal2 s 57792 59600 57848 59900 6 io_in[12]
port 4 nsew signal input
rlabel metal3 s 100 21168 400 21224 6 io_in[13]
port 5 nsew signal input
rlabel metal2 s 32928 59600 32984 59900 6 io_in[14]
port 6 nsew signal input
rlabel metal3 s 59600 11424 59900 11480 6 io_in[15]
port 7 nsew signal input
rlabel metal2 s 17136 100 17192 400 6 io_in[16]
port 8 nsew signal input
rlabel metal2 s 13440 59600 13496 59900 6 io_in[17]
port 9 nsew signal input
rlabel metal3 s 100 26544 400 26600 6 io_in[18]
port 10 nsew signal input
rlabel metal3 s 59600 59808 59900 59864 6 io_in[19]
port 11 nsew signal input
rlabel metal2 s 48048 59600 48104 59900 6 io_in[1]
port 12 nsew signal input
rlabel metal2 s 34608 59600 34664 59900 6 io_in[20]
port 13 nsew signal input
rlabel metal2 s 56784 59600 56840 59900 6 io_in[21]
port 14 nsew signal input
rlabel metal2 s 1008 59600 1064 59900 6 io_in[22]
port 15 nsew signal input
rlabel metal2 s 8064 100 8120 400 6 io_in[23]
port 16 nsew signal input
rlabel metal2 s 7392 59600 7448 59900 6 io_in[24]
port 17 nsew signal input
rlabel metal2 s 9744 59600 9800 59900 6 io_in[25]
port 18 nsew signal input
rlabel metal3 s 59600 6384 59900 6440 6 io_in[26]
port 19 nsew signal input
rlabel metal3 s 100 14448 400 14504 6 io_in[27]
port 20 nsew signal input
rlabel metal2 s 2352 59600 2408 59900 6 io_in[28]
port 21 nsew signal input
rlabel metal3 s 59600 58464 59900 58520 6 io_in[29]
port 22 nsew signal input
rlabel metal3 s 100 6048 400 6104 6 io_in[2]
port 23 nsew signal input
rlabel metal2 s 42000 100 42056 400 6 io_in[30]
port 24 nsew signal input
rlabel metal2 s 8736 59600 8792 59900 6 io_in[31]
port 25 nsew signal input
rlabel metal2 s 35616 100 35672 400 6 io_in[32]
port 26 nsew signal input
rlabel metal3 s 100 58800 400 58856 6 io_in[33]
port 27 nsew signal input
rlabel metal2 s 53760 59600 53816 59900 6 io_in[34]
port 28 nsew signal input
rlabel metal2 s 12768 59600 12824 59900 6 io_in[35]
port 29 nsew signal input
rlabel metal3 s 100 15456 400 15512 6 io_in[36]
port 30 nsew signal input
rlabel metal3 s 59600 9744 59900 9800 6 io_in[37]
port 31 nsew signal input
rlabel metal3 s 100 25200 400 25256 6 io_in[3]
port 32 nsew signal input
rlabel metal2 s 53760 100 53816 400 6 io_in[4]
port 33 nsew signal input
rlabel metal3 s 100 58464 400 58520 6 io_in[5]
port 34 nsew signal input
rlabel metal3 s 100 13776 400 13832 6 io_in[6]
port 35 nsew signal input
rlabel metal3 s 59600 15792 59900 15848 6 io_in[7]
port 36 nsew signal input
rlabel metal2 s 58464 100 58520 400 6 io_in[8]
port 37 nsew signal input
rlabel metal2 s 51072 59600 51128 59900 6 io_in[9]
port 38 nsew signal input
rlabel metal2 s 1680 59600 1736 59900 6 io_oeb[0]
port 39 nsew signal output
rlabel metal3 s 100 40992 400 41048 6 io_oeb[10]
port 40 nsew signal output
rlabel metal3 s 100 37632 400 37688 6 io_oeb[11]
port 41 nsew signal output
rlabel metal3 s 100 45024 400 45080 6 io_oeb[12]
port 42 nsew signal output
rlabel metal2 s 51408 100 51464 400 6 io_oeb[13]
port 43 nsew signal output
rlabel metal2 s 58800 100 58856 400 6 io_oeb[14]
port 44 nsew signal output
rlabel metal2 s 31920 59600 31976 59900 6 io_oeb[15]
port 45 nsew signal output
rlabel metal3 s 100 34608 400 34664 6 io_oeb[16]
port 46 nsew signal output
rlabel metal2 s 5712 59600 5768 59900 6 io_oeb[17]
port 47 nsew signal output
rlabel metal3 s 100 47376 400 47432 6 io_oeb[18]
port 48 nsew signal output
rlabel metal2 s 24192 100 24248 400 6 io_oeb[19]
port 49 nsew signal output
rlabel metal3 s 59600 4704 59900 4760 6 io_oeb[1]
port 50 nsew signal output
rlabel metal2 s 50736 100 50792 400 6 io_oeb[20]
port 51 nsew signal output
rlabel metal2 s 5712 100 5768 400 6 io_oeb[21]
port 52 nsew signal output
rlabel metal3 s 59600 15120 59900 15176 6 io_oeb[22]
port 53 nsew signal output
rlabel metal3 s 100 5712 400 5768 6 io_oeb[23]
port 54 nsew signal output
rlabel metal3 s 59600 13440 59900 13496 6 io_oeb[24]
port 55 nsew signal output
rlabel metal2 s 21168 100 21224 400 6 io_oeb[25]
port 56 nsew signal output
rlabel metal2 s 49728 100 49784 400 6 io_oeb[26]
port 57 nsew signal output
rlabel metal3 s 100 39984 400 40040 6 io_oeb[27]
port 58 nsew signal output
rlabel metal3 s 100 56112 400 56168 6 io_oeb[28]
port 59 nsew signal output
rlabel metal2 s 12096 59600 12152 59900 6 io_oeb[29]
port 60 nsew signal output
rlabel metal2 s 38640 100 38696 400 6 io_oeb[2]
port 61 nsew signal output
rlabel metal3 s 100 2016 400 2072 6 io_oeb[30]
port 62 nsew signal output
rlabel metal3 s 59600 41664 59900 41720 6 io_oeb[31]
port 63 nsew signal output
rlabel metal3 s 59600 9408 59900 9464 6 io_oeb[32]
port 64 nsew signal output
rlabel metal3 s 100 49056 400 49112 6 io_oeb[33]
port 65 nsew signal output
rlabel metal3 s 100 23184 400 23240 6 io_oeb[34]
port 66 nsew signal output
rlabel metal2 s 33600 59600 33656 59900 6 io_oeb[35]
port 67 nsew signal output
rlabel metal2 s 56112 100 56168 400 6 io_oeb[36]
port 68 nsew signal output
rlabel metal3 s 100 50400 400 50456 6 io_oeb[37]
port 69 nsew signal output
rlabel metal3 s 59600 20160 59900 20216 6 io_oeb[3]
port 70 nsew signal output
rlabel metal2 s 0 59600 56 59900 6 io_oeb[4]
port 71 nsew signal output
rlabel metal3 s 59600 57792 59900 57848 6 io_oeb[5]
port 72 nsew signal output
rlabel metal2 s 28896 59600 28952 59900 6 io_oeb[6]
port 73 nsew signal output
rlabel metal3 s 59600 3360 59900 3416 6 io_oeb[7]
port 74 nsew signal output
rlabel metal3 s 59600 24192 59900 24248 6 io_oeb[8]
port 75 nsew signal output
rlabel metal3 s 59600 23856 59900 23912 6 io_oeb[9]
port 76 nsew signal output
rlabel metal3 s 100 11424 400 11480 6 io_out[0]
port 77 nsew signal output
rlabel metal2 s 58464 59600 58520 59900 6 io_out[10]
port 78 nsew signal output
rlabel metal3 s 59600 52752 59900 52808 6 io_out[11]
port 79 nsew signal output
rlabel metal3 s 59600 59136 59900 59192 6 io_out[12]
port 80 nsew signal output
rlabel metal3 s 100 44352 400 44408 6 io_out[13]
port 81 nsew signal output
rlabel metal2 s 23520 100 23576 400 6 io_out[14]
port 82 nsew signal output
rlabel metal3 s 59600 49728 59900 49784 6 io_out[15]
port 83 nsew signal output
rlabel metal2 s 6720 100 6776 400 6 io_out[16]
port 84 nsew signal output
rlabel metal2 s 50400 100 50456 400 6 io_out[17]
port 85 nsew signal output
rlabel metal2 s 39312 100 39368 400 6 io_out[18]
port 86 nsew signal output
rlabel metal2 s 4032 100 4088 400 6 io_out[19]
port 87 nsew signal output
rlabel metal2 s 40992 100 41048 400 6 io_out[1]
port 88 nsew signal output
rlabel metal2 s 27216 100 27272 400 6 io_out[20]
port 89 nsew signal output
rlabel metal2 s 20160 100 20216 400 6 io_out[21]
port 90 nsew signal output
rlabel metal3 s 100 8064 400 8120 6 io_out[22]
port 91 nsew signal output
rlabel metal2 s 44016 59600 44072 59900 6 io_out[23]
port 92 nsew signal output
rlabel metal2 s 27888 59600 27944 59900 6 io_out[24]
port 93 nsew signal output
rlabel metal2 s 25200 100 25256 400 6 io_out[25]
port 94 nsew signal output
rlabel metal2 s 42336 59600 42392 59900 6 io_out[26]
port 95 nsew signal output
rlabel metal2 s 44352 100 44408 400 6 io_out[27]
port 96 nsew signal output
rlabel metal2 s 38304 59600 38360 59900 6 io_out[28]
port 97 nsew signal output
rlabel metal2 s 56784 100 56840 400 6 io_out[29]
port 98 nsew signal output
rlabel metal2 s 55104 59600 55160 59900 6 io_out[2]
port 99 nsew signal output
rlabel metal3 s 59600 12768 59900 12824 6 io_out[30]
port 100 nsew signal output
rlabel metal2 s 50400 59600 50456 59900 6 io_out[31]
port 101 nsew signal output
rlabel metal3 s 59600 19152 59900 19208 6 io_out[32]
port 102 nsew signal output
rlabel metal2 s 39984 100 40040 400 6 io_out[33]
port 103 nsew signal output
rlabel metal3 s 59600 38976 59900 39032 6 io_out[34]
port 104 nsew signal output
rlabel metal2 s 14448 100 14504 400 6 io_out[35]
port 105 nsew signal output
rlabel metal3 s 59600 56112 59900 56168 6 io_out[36]
port 106 nsew signal output
rlabel metal3 s 59600 55776 59900 55832 6 io_out[37]
port 107 nsew signal output
rlabel metal3 s 59600 43008 59900 43064 6 io_out[3]
port 108 nsew signal output
rlabel metal3 s 100 1680 400 1736 6 io_out[4]
port 109 nsew signal output
rlabel metal3 s 100 2688 400 2744 6 io_out[5]
port 110 nsew signal output
rlabel metal3 s 100 33936 400 33992 6 io_out[6]
port 111 nsew signal output
rlabel metal2 s 37632 59600 37688 59900 6 io_out[7]
port 112 nsew signal output
rlabel metal2 s 15456 100 15512 400 6 io_out[8]
port 113 nsew signal output
rlabel metal3 s 100 30576 400 30632 6 io_out[9]
port 114 nsew signal output
rlabel metal3 s 100 42000 400 42056 6 irq[0]
port 115 nsew signal output
rlabel metal3 s 100 24192 400 24248 6 irq[1]
port 116 nsew signal output
rlabel metal2 s 18480 100 18536 400 6 irq[2]
port 117 nsew signal output
rlabel metal2 s 24192 59600 24248 59900 6 la_data_in[0]
port 118 nsew signal input
rlabel metal2 s 56112 59600 56168 59900 6 la_data_in[10]
port 119 nsew signal input
rlabel metal2 s 28224 100 28280 400 6 la_data_in[11]
port 120 nsew signal input
rlabel metal3 s 100 36288 400 36344 6 la_data_in[12]
port 121 nsew signal input
rlabel metal3 s 59600 8736 59900 8792 6 la_data_in[13]
port 122 nsew signal input
rlabel metal3 s 59600 21840 59900 21896 6 la_data_in[14]
port 123 nsew signal input
rlabel metal3 s 100 41664 400 41720 6 la_data_in[15]
port 124 nsew signal input
rlabel metal2 s 13776 59600 13832 59900 6 la_data_in[16]
port 125 nsew signal input
rlabel metal3 s 59600 12096 59900 12152 6 la_data_in[17]
port 126 nsew signal input
rlabel metal3 s 59600 45360 59900 45416 6 la_data_in[18]
port 127 nsew signal input
rlabel metal3 s 59600 26544 59900 26600 6 la_data_in[19]
port 128 nsew signal input
rlabel metal2 s 45696 59600 45752 59900 6 la_data_in[1]
port 129 nsew signal input
rlabel metal2 s 30576 59600 30632 59900 6 la_data_in[20]
port 130 nsew signal input
rlabel metal3 s 100 9744 400 9800 6 la_data_in[21]
port 131 nsew signal input
rlabel metal2 s 36960 59600 37016 59900 6 la_data_in[22]
port 132 nsew signal input
rlabel metal3 s 100 54432 400 54488 6 la_data_in[23]
port 133 nsew signal input
rlabel metal2 s 26208 59600 26264 59900 6 la_data_in[24]
port 134 nsew signal input
rlabel metal3 s 59600 14448 59900 14504 6 la_data_in[25]
port 135 nsew signal input
rlabel metal2 s 19488 100 19544 400 6 la_data_in[26]
port 136 nsew signal input
rlabel metal3 s 100 4368 400 4424 6 la_data_in[27]
port 137 nsew signal input
rlabel metal3 s 100 21840 400 21896 6 la_data_in[28]
port 138 nsew signal input
rlabel metal3 s 100 45696 400 45752 6 la_data_in[29]
port 139 nsew signal input
rlabel metal3 s 100 40320 400 40376 6 la_data_in[2]
port 140 nsew signal input
rlabel metal2 s 4704 59600 4760 59900 6 la_data_in[30]
port 141 nsew signal input
rlabel metal3 s 100 53088 400 53144 6 la_data_in[31]
port 142 nsew signal input
rlabel metal2 s 30240 59600 30296 59900 6 la_data_in[32]
port 143 nsew signal input
rlabel metal3 s 59600 51072 59900 51128 6 la_data_in[33]
port 144 nsew signal input
rlabel metal2 s 18480 59600 18536 59900 6 la_data_in[34]
port 145 nsew signal input
rlabel metal2 s 24864 59600 24920 59900 6 la_data_in[35]
port 146 nsew signal input
rlabel metal3 s 59600 32592 59900 32648 6 la_data_in[36]
port 147 nsew signal input
rlabel metal2 s 20832 100 20888 400 6 la_data_in[37]
port 148 nsew signal input
rlabel metal2 s 28896 100 28952 400 6 la_data_in[38]
port 149 nsew signal input
rlabel metal3 s 100 20160 400 20216 6 la_data_in[39]
port 150 nsew signal input
rlabel metal3 s 59600 36960 59900 37016 6 la_data_in[3]
port 151 nsew signal input
rlabel metal3 s 59600 672 59900 728 6 la_data_in[40]
port 152 nsew signal input
rlabel metal3 s 100 56784 400 56840 6 la_data_in[41]
port 153 nsew signal input
rlabel metal3 s 59600 43344 59900 43400 6 la_data_in[42]
port 154 nsew signal input
rlabel metal2 s 36960 100 37016 400 6 la_data_in[43]
port 155 nsew signal input
rlabel metal2 s 28224 59600 28280 59900 6 la_data_in[44]
port 156 nsew signal input
rlabel metal2 s 8064 59600 8120 59900 6 la_data_in[45]
port 157 nsew signal input
rlabel metal2 s 5040 59600 5096 59900 6 la_data_in[46]
port 158 nsew signal input
rlabel metal2 s 23856 59600 23912 59900 6 la_data_in[47]
port 159 nsew signal input
rlabel metal2 s 27552 100 27608 400 6 la_data_in[48]
port 160 nsew signal input
rlabel metal3 s 100 31248 400 31304 6 la_data_in[49]
port 161 nsew signal input
rlabel metal2 s 49392 59600 49448 59900 6 la_data_in[4]
port 162 nsew signal input
rlabel metal3 s 100 18480 400 18536 6 la_data_in[50]
port 163 nsew signal input
rlabel metal3 s 100 16128 400 16184 6 la_data_in[51]
port 164 nsew signal input
rlabel metal3 s 100 17808 400 17864 6 la_data_in[52]
port 165 nsew signal input
rlabel metal3 s 59600 1680 59900 1736 6 la_data_in[53]
port 166 nsew signal input
rlabel metal2 s 21840 100 21896 400 6 la_data_in[54]
port 167 nsew signal input
rlabel metal3 s 59600 54432 59900 54488 6 la_data_in[55]
port 168 nsew signal input
rlabel metal2 s 10416 100 10472 400 6 la_data_in[56]
port 169 nsew signal input
rlabel metal2 s 15792 59600 15848 59900 6 la_data_in[57]
port 170 nsew signal input
rlabel metal2 s 22512 59600 22568 59900 6 la_data_in[58]
port 171 nsew signal input
rlabel metal2 s 35280 100 35336 400 6 la_data_in[59]
port 172 nsew signal input
rlabel metal3 s 100 336 400 392 6 la_data_in[5]
port 173 nsew signal input
rlabel metal2 s 12096 100 12152 400 6 la_data_in[60]
port 174 nsew signal input
rlabel metal3 s 59600 21504 59900 21560 6 la_data_in[61]
port 175 nsew signal input
rlabel metal2 s 17808 59600 17864 59900 6 la_data_in[62]
port 176 nsew signal input
rlabel metal2 s 54432 59600 54488 59900 6 la_data_in[63]
port 177 nsew signal input
rlabel metal2 s 52080 59600 52136 59900 6 la_data_in[6]
port 178 nsew signal input
rlabel metal3 s 59600 31920 59900 31976 6 la_data_in[7]
port 179 nsew signal input
rlabel metal2 s 42672 100 42728 400 6 la_data_in[8]
port 180 nsew signal input
rlabel metal3 s 100 43344 400 43400 6 la_data_in[9]
port 181 nsew signal input
rlabel metal2 s 16800 59600 16856 59900 6 la_data_out[0]
port 182 nsew signal output
rlabel metal3 s 59600 24864 59900 24920 6 la_data_out[10]
port 183 nsew signal output
rlabel metal3 s 100 51408 400 51464 6 la_data_out[11]
port 184 nsew signal output
rlabel metal3 s 59600 32928 59900 32984 6 la_data_out[12]
port 185 nsew signal output
rlabel metal2 s 29568 59600 29624 59900 6 la_data_out[13]
port 186 nsew signal output
rlabel metal2 s 26544 59600 26600 59900 6 la_data_out[14]
port 187 nsew signal output
rlabel metal2 s 31584 100 31640 400 6 la_data_out[15]
port 188 nsew signal output
rlabel metal3 s 59600 27888 59900 27944 6 la_data_out[16]
port 189 nsew signal output
rlabel metal2 s 59136 59600 59192 59900 6 la_data_out[17]
port 190 nsew signal output
rlabel metal3 s 100 59472 400 59528 6 la_data_out[18]
port 191 nsew signal output
rlabel metal3 s 59600 37632 59900 37688 6 la_data_out[19]
port 192 nsew signal output
rlabel metal2 s 17808 100 17864 400 6 la_data_out[1]
port 193 nsew signal output
rlabel metal3 s 59600 17472 59900 17528 6 la_data_out[20]
port 194 nsew signal output
rlabel metal3 s 100 10416 400 10472 6 la_data_out[21]
port 195 nsew signal output
rlabel metal3 s 59600 7392 59900 7448 6 la_data_out[22]
port 196 nsew signal output
rlabel metal2 s 36624 59600 36680 59900 6 la_data_out[23]
port 197 nsew signal output
rlabel metal3 s 59600 47376 59900 47432 6 la_data_out[24]
port 198 nsew signal output
rlabel metal2 s 25872 100 25928 400 6 la_data_out[25]
port 199 nsew signal output
rlabel metal3 s 100 46704 400 46760 6 la_data_out[26]
port 200 nsew signal output
rlabel metal3 s 59600 27216 59900 27272 6 la_data_out[27]
port 201 nsew signal output
rlabel metal3 s 100 22512 400 22568 6 la_data_out[28]
port 202 nsew signal output
rlabel metal2 s 35280 59600 35336 59900 6 la_data_out[29]
port 203 nsew signal output
rlabel metal3 s 59600 11088 59900 11144 6 la_data_out[2]
port 204 nsew signal output
rlabel metal2 s 29232 100 29288 400 6 la_data_out[30]
port 205 nsew signal output
rlabel metal2 s 32592 59600 32648 59900 6 la_data_out[31]
port 206 nsew signal output
rlabel metal3 s 59600 48048 59900 48104 6 la_data_out[32]
port 207 nsew signal output
rlabel metal3 s 59600 23184 59900 23240 6 la_data_out[33]
port 208 nsew signal output
rlabel metal3 s 59600 1008 59900 1064 6 la_data_out[34]
port 209 nsew signal output
rlabel metal3 s 59600 8064 59900 8120 6 la_data_out[35]
port 210 nsew signal output
rlabel metal3 s 100 3360 400 3416 6 la_data_out[36]
port 211 nsew signal output
rlabel metal3 s 100 53760 400 53816 6 la_data_out[37]
port 212 nsew signal output
rlabel metal3 s 100 27216 400 27272 6 la_data_out[38]
port 213 nsew signal output
rlabel metal3 s 59600 50400 59900 50456 6 la_data_out[39]
port 214 nsew signal output
rlabel metal2 s 3360 100 3416 400 6 la_data_out[3]
port 215 nsew signal output
rlabel metal2 s 24864 100 24920 400 6 la_data_out[40]
port 216 nsew signal output
rlabel metal2 s 9408 59600 9464 59900 6 la_data_out[41]
port 217 nsew signal output
rlabel metal2 s 54768 100 54824 400 6 la_data_out[42]
port 218 nsew signal output
rlabel metal3 s 100 42672 400 42728 6 la_data_out[43]
port 219 nsew signal output
rlabel metal2 s 13776 100 13832 400 6 la_data_out[44]
port 220 nsew signal output
rlabel metal2 s 54432 100 54488 400 6 la_data_out[45]
port 221 nsew signal output
rlabel metal2 s 34272 59600 34328 59900 6 la_data_out[46]
port 222 nsew signal output
rlabel metal2 s 20832 59600 20888 59900 6 la_data_out[47]
port 223 nsew signal output
rlabel metal3 s 100 57792 400 57848 6 la_data_out[48]
port 224 nsew signal output
rlabel metal2 s 43344 59600 43400 59900 6 la_data_out[49]
port 225 nsew signal output
rlabel metal3 s 100 1008 400 1064 6 la_data_out[4]
port 226 nsew signal output
rlabel metal2 s 47040 59600 47096 59900 6 la_data_out[50]
port 227 nsew signal output
rlabel metal2 s 25536 59600 25592 59900 6 la_data_out[51]
port 228 nsew signal output
rlabel metal3 s 100 8400 400 8456 6 la_data_out[52]
port 229 nsew signal output
rlabel metal3 s 59600 35280 59900 35336 6 la_data_out[53]
port 230 nsew signal output
rlabel metal3 s 59600 40992 59900 41048 6 la_data_out[54]
port 231 nsew signal output
rlabel metal3 s 59600 53424 59900 53480 6 la_data_out[55]
port 232 nsew signal output
rlabel metal3 s 100 54768 400 54824 6 la_data_out[56]
port 233 nsew signal output
rlabel metal2 s 48720 59600 48776 59900 6 la_data_out[57]
port 234 nsew signal output
rlabel metal2 s 16128 100 16184 400 6 la_data_out[58]
port 235 nsew signal output
rlabel metal2 s 52080 100 52136 400 6 la_data_out[59]
port 236 nsew signal output
rlabel metal3 s 59600 4032 59900 4088 6 la_data_out[5]
port 237 nsew signal output
rlabel metal3 s 100 9072 400 9128 6 la_data_out[60]
port 238 nsew signal output
rlabel metal2 s 21504 59600 21560 59900 6 la_data_out[61]
port 239 nsew signal output
rlabel metal2 s 37632 100 37688 400 6 la_data_out[62]
port 240 nsew signal output
rlabel metal3 s 59600 28224 59900 28280 6 la_data_out[63]
port 241 nsew signal output
rlabel metal3 s 59600 22512 59900 22568 6 la_data_out[6]
port 242 nsew signal output
rlabel metal3 s 59600 42336 59900 42392 6 la_data_out[7]
port 243 nsew signal output
rlabel metal3 s 59600 33600 59900 33656 6 la_data_out[8]
port 244 nsew signal output
rlabel metal2 s 23184 59600 23240 59900 6 la_data_out[9]
port 245 nsew signal output
rlabel metal3 s 100 48048 400 48104 6 la_oenb[0]
port 246 nsew signal input
rlabel metal2 s 44016 100 44072 400 6 la_oenb[10]
port 247 nsew signal input
rlabel metal2 s 52752 100 52808 400 6 la_oenb[11]
port 248 nsew signal input
rlabel metal2 s 8400 100 8456 400 6 la_oenb[12]
port 249 nsew signal input
rlabel metal3 s 100 7392 400 7448 6 la_oenb[13]
port 250 nsew signal input
rlabel metal2 s 4032 59600 4088 59900 6 la_oenb[14]
port 251 nsew signal input
rlabel metal3 s 59600 5040 59900 5096 6 la_oenb[15]
port 252 nsew signal input
rlabel metal2 s 11424 59600 11480 59900 6 la_oenb[16]
port 253 nsew signal input
rlabel metal3 s 100 52752 400 52808 6 la_oenb[17]
port 254 nsew signal input
rlabel metal2 s 52752 59600 52808 59900 6 la_oenb[18]
port 255 nsew signal input
rlabel metal2 s 44688 59600 44744 59900 6 la_oenb[19]
port 256 nsew signal input
rlabel metal2 s 16800 100 16856 400 6 la_oenb[1]
port 257 nsew signal input
rlabel metal3 s 100 33600 400 33656 6 la_oenb[20]
port 258 nsew signal input
rlabel metal2 s 53088 100 53144 400 6 la_oenb[21]
port 259 nsew signal input
rlabel metal3 s 100 32256 400 32312 6 la_oenb[22]
port 260 nsew signal input
rlabel metal2 s 10752 100 10808 400 6 la_oenb[23]
port 261 nsew signal input
rlabel metal3 s 100 36960 400 37016 6 la_oenb[24]
port 262 nsew signal input
rlabel metal3 s 59600 56784 59900 56840 6 la_oenb[25]
port 263 nsew signal input
rlabel metal2 s 59808 59600 59864 59900 6 la_oenb[26]
port 264 nsew signal input
rlabel metal3 s 59600 51408 59900 51464 6 la_oenb[27]
port 265 nsew signal input
rlabel metal3 s 59600 49392 59900 49448 6 la_oenb[28]
port 266 nsew signal input
rlabel metal3 s 59600 48720 59900 48776 6 la_oenb[29]
port 267 nsew signal input
rlabel metal2 s 30576 100 30632 400 6 la_oenb[2]
port 268 nsew signal input
rlabel metal2 s 10416 59600 10472 59900 6 la_oenb[30]
port 269 nsew signal input
rlabel metal2 s 1680 100 1736 400 6 la_oenb[31]
port 270 nsew signal input
rlabel metal2 s 336 100 392 400 6 la_oenb[32]
port 271 nsew signal input
rlabel metal2 s 672 59600 728 59900 6 la_oenb[33]
port 272 nsew signal input
rlabel metal2 s 31248 100 31304 400 6 la_oenb[34]
port 273 nsew signal input
rlabel metal3 s 100 25872 400 25928 6 la_oenb[35]
port 274 nsew signal input
rlabel metal3 s 100 32928 400 32984 6 la_oenb[36]
port 275 nsew signal input
rlabel metal3 s 100 17136 400 17192 6 la_oenb[37]
port 276 nsew signal input
rlabel metal2 s 21840 59600 21896 59900 6 la_oenb[38]
port 277 nsew signal input
rlabel metal3 s 100 37968 400 38024 6 la_oenb[39]
port 278 nsew signal input
rlabel metal2 s 11424 100 11480 400 6 la_oenb[3]
port 279 nsew signal input
rlabel metal2 s 26544 100 26600 400 6 la_oenb[40]
port 280 nsew signal input
rlabel metal3 s 100 29904 400 29960 6 la_oenb[41]
port 281 nsew signal input
rlabel metal2 s 48048 100 48104 400 6 la_oenb[42]
port 282 nsew signal input
rlabel metal2 s 22512 100 22568 400 6 la_oenb[43]
port 283 nsew signal input
rlabel metal3 s 100 44016 400 44072 6 la_oenb[44]
port 284 nsew signal input
rlabel metal3 s 59600 28896 59900 28952 6 la_oenb[45]
port 285 nsew signal input
rlabel metal3 s 59600 39984 59900 40040 6 la_oenb[46]
port 286 nsew signal input
rlabel metal2 s 46368 100 46424 400 6 la_oenb[47]
port 287 nsew signal input
rlabel metal2 s 19824 59600 19880 59900 6 la_oenb[48]
port 288 nsew signal input
rlabel metal2 s 59472 100 59528 400 6 la_oenb[49]
port 289 nsew signal input
rlabel metal3 s 59600 38304 59900 38360 6 la_oenb[4]
port 290 nsew signal input
rlabel metal2 s 40656 59600 40712 59900 6 la_oenb[50]
port 291 nsew signal input
rlabel metal3 s 59600 30576 59900 30632 6 la_oenb[51]
port 292 nsew signal input
rlabel metal2 s 45696 100 45752 400 6 la_oenb[52]
port 293 nsew signal input
rlabel metal2 s 53424 59600 53480 59900 6 la_oenb[53]
port 294 nsew signal input
rlabel metal3 s 59600 5712 59900 5768 6 la_oenb[54]
port 295 nsew signal input
rlabel metal2 s 35952 59600 36008 59900 6 la_oenb[55]
port 296 nsew signal input
rlabel metal2 s 55440 100 55496 400 6 la_oenb[56]
port 297 nsew signal input
rlabel metal3 s 100 29232 400 29288 6 la_oenb[57]
port 298 nsew signal input
rlabel metal2 s 7392 100 7448 400 6 la_oenb[58]
port 299 nsew signal input
rlabel metal3 s 59600 30240 59900 30296 6 la_oenb[59]
port 300 nsew signal input
rlabel metal3 s 100 57120 400 57176 6 la_oenb[5]
port 301 nsew signal input
rlabel metal3 s 59600 39312 59900 39368 6 la_oenb[60]
port 302 nsew signal input
rlabel metal2 s 14784 100 14840 400 6 la_oenb[61]
port 303 nsew signal input
rlabel metal2 s 57120 100 57176 400 6 la_oenb[62]
port 304 nsew signal input
rlabel metal3 s 100 10752 400 10808 6 la_oenb[63]
port 305 nsew signal input
rlabel metal2 s 51408 59600 51464 59900 6 la_oenb[6]
port 306 nsew signal input
rlabel metal3 s 59600 45696 59900 45752 6 la_oenb[7]
port 307 nsew signal input
rlabel metal2 s 15120 59600 15176 59900 6 la_oenb[8]
port 308 nsew signal input
rlabel metal3 s 100 38640 400 38696 6 la_oenb[9]
port 309 nsew signal input
rlabel metal4 s 2224 1538 2384 58438 6 vdd
port 310 nsew power bidirectional
rlabel metal4 s 17584 1538 17744 58438 6 vdd
port 310 nsew power bidirectional
rlabel metal4 s 32944 1538 33104 58438 6 vdd
port 310 nsew power bidirectional
rlabel metal4 s 48304 1538 48464 58438 6 vdd
port 310 nsew power bidirectional
rlabel metal4 s 9904 1538 10064 58438 6 vss
port 311 nsew ground bidirectional
rlabel metal4 s 25264 1538 25424 58438 6 vss
port 311 nsew ground bidirectional
rlabel metal4 s 40624 1538 40784 58438 6 vss
port 311 nsew ground bidirectional
rlabel metal4 s 55984 1538 56144 58438 6 vss
port 311 nsew ground bidirectional
rlabel metal3 s 59600 10416 59900 10472 6 wb_clk_i
port 312 nsew signal input
rlabel metal2 s 11088 59600 11144 59900 6 wb_rst_i
port 313 nsew signal input
rlabel metal3 s 59600 20832 59900 20888 6 wbs_ack_o
port 314 nsew signal output
rlabel metal2 s 39984 59600 40040 59900 6 wbs_adr_i[0]
port 315 nsew signal input
rlabel metal2 s 27216 59600 27272 59900 6 wbs_adr_i[10]
port 316 nsew signal input
rlabel metal2 s 3360 59600 3416 59900 6 wbs_adr_i[11]
port 317 nsew signal input
rlabel metal2 s 5040 100 5096 400 6 wbs_adr_i[12]
port 318 nsew signal input
rlabel metal2 s 33600 100 33656 400 6 wbs_adr_i[13]
port 319 nsew signal input
rlabel metal3 s 59600 44016 59900 44072 6 wbs_adr_i[14]
port 320 nsew signal input
rlabel metal3 s 59600 40656 59900 40712 6 wbs_adr_i[15]
port 321 nsew signal input
rlabel metal2 s 37968 100 38024 400 6 wbs_adr_i[16]
port 322 nsew signal input
rlabel metal3 s 59600 35952 59900 36008 6 wbs_adr_i[17]
port 323 nsew signal input
rlabel metal3 s 59600 18480 59900 18536 6 wbs_adr_i[18]
port 324 nsew signal input
rlabel metal2 s 57792 100 57848 400 6 wbs_adr_i[19]
port 325 nsew signal input
rlabel metal3 s 100 4032 400 4088 6 wbs_adr_i[1]
port 326 nsew signal input
rlabel metal3 s 100 35280 400 35336 6 wbs_adr_i[20]
port 327 nsew signal input
rlabel metal2 s 33936 100 33992 400 6 wbs_adr_i[21]
port 328 nsew signal input
rlabel metal2 s 48384 100 48440 400 6 wbs_adr_i[22]
port 329 nsew signal input
rlabel metal3 s 59600 13776 59900 13832 6 wbs_adr_i[23]
port 330 nsew signal input
rlabel metal2 s 7056 59600 7112 59900 6 wbs_adr_i[24]
port 331 nsew signal input
rlabel metal2 s 32928 100 32984 400 6 wbs_adr_i[25]
port 332 nsew signal input
rlabel metal2 s 6048 100 6104 400 6 wbs_adr_i[26]
port 333 nsew signal input
rlabel metal2 s 20160 59600 20216 59900 6 wbs_adr_i[27]
port 334 nsew signal input
rlabel metal3 s 59600 34608 59900 34664 6 wbs_adr_i[28]
port 335 nsew signal input
rlabel metal3 s 59600 57456 59900 57512 6 wbs_adr_i[29]
port 336 nsew signal input
rlabel metal3 s 100 6720 400 6776 6 wbs_adr_i[2]
port 337 nsew signal input
rlabel metal3 s 100 23520 400 23576 6 wbs_adr_i[30]
port 338 nsew signal input
rlabel metal3 s 59600 25536 59900 25592 6 wbs_adr_i[31]
port 339 nsew signal input
rlabel metal2 s 46704 100 46760 400 6 wbs_adr_i[3]
port 340 nsew signal input
rlabel metal2 s 46368 59600 46424 59900 6 wbs_adr_i[4]
port 341 nsew signal input
rlabel metal2 s 45024 100 45080 400 6 wbs_adr_i[5]
port 342 nsew signal input
rlabel metal3 s 100 28896 400 28952 6 wbs_adr_i[6]
port 343 nsew signal input
rlabel metal2 s 2688 100 2744 400 6 wbs_adr_i[7]
port 344 nsew signal input
rlabel metal3 s 59600 0 59900 56 6 wbs_adr_i[8]
port 345 nsew signal input
rlabel metal3 s 59600 16128 59900 16184 6 wbs_adr_i[9]
port 346 nsew signal input
rlabel metal2 s 19152 59600 19208 59900 6 wbs_cyc_i
port 347 nsew signal input
rlabel metal3 s 59600 52080 59900 52136 6 wbs_dat_i[0]
port 348 nsew signal input
rlabel metal3 s 100 46368 400 46424 6 wbs_dat_i[10]
port 349 nsew signal input
rlabel metal3 s 100 50736 400 50792 6 wbs_dat_i[11]
port 350 nsew signal input
rlabel metal3 s 100 48384 400 48440 6 wbs_dat_i[12]
port 351 nsew signal input
rlabel metal2 s 2016 100 2072 400 6 wbs_dat_i[13]
port 352 nsew signal input
rlabel metal3 s 100 12432 400 12488 6 wbs_dat_i[14]
port 353 nsew signal input
rlabel metal3 s 59600 31248 59900 31304 6 wbs_dat_i[15]
port 354 nsew signal input
rlabel metal2 s 34608 100 34664 400 6 wbs_dat_i[16]
port 355 nsew signal input
rlabel metal2 s 40992 59600 41048 59900 6 wbs_dat_i[17]
port 356 nsew signal input
rlabel metal2 s 55776 59600 55832 59900 6 wbs_dat_i[18]
port 357 nsew signal input
rlabel metal2 s 3024 59600 3080 59900 6 wbs_dat_i[19]
port 358 nsew signal input
rlabel metal2 s 9072 100 9128 400 6 wbs_dat_i[1]
port 359 nsew signal input
rlabel metal3 s 100 14784 400 14840 6 wbs_dat_i[20]
port 360 nsew signal input
rlabel metal2 s 57456 59600 57512 59900 6 wbs_dat_i[21]
port 361 nsew signal input
rlabel metal3 s 100 35616 400 35672 6 wbs_dat_i[22]
port 362 nsew signal input
rlabel metal3 s 59600 47040 59900 47096 6 wbs_dat_i[23]
port 363 nsew signal input
rlabel metal3 s 59600 19824 59900 19880 6 wbs_dat_i[24]
port 364 nsew signal input
rlabel metal2 s 41664 100 41720 400 6 wbs_dat_i[25]
port 365 nsew signal input
rlabel metal2 s 49728 59600 49784 59900 6 wbs_dat_i[26]
port 366 nsew signal input
rlabel metal2 s 14448 59600 14504 59900 6 wbs_dat_i[27]
port 367 nsew signal input
rlabel metal2 s 18816 100 18872 400 6 wbs_dat_i[28]
port 368 nsew signal input
rlabel metal3 s 59600 36624 59900 36680 6 wbs_dat_i[29]
port 369 nsew signal input
rlabel metal2 s 49056 100 49112 400 6 wbs_dat_i[2]
port 370 nsew signal input
rlabel metal3 s 59600 17808 59900 17864 6 wbs_dat_i[30]
port 371 nsew signal input
rlabel metal3 s 100 31584 400 31640 6 wbs_dat_i[31]
port 372 nsew signal input
rlabel metal3 s 59600 2352 59900 2408 6 wbs_dat_i[3]
port 373 nsew signal input
rlabel metal2 s 9744 100 9800 400 6 wbs_dat_i[4]
port 374 nsew signal input
rlabel metal2 s 29904 100 29960 400 6 wbs_dat_i[5]
port 375 nsew signal input
rlabel metal3 s 59600 26208 59900 26264 6 wbs_dat_i[6]
port 376 nsew signal input
rlabel metal2 s 47376 59600 47432 59900 6 wbs_dat_i[7]
port 377 nsew signal input
rlabel metal3 s 59600 53760 59900 53816 6 wbs_dat_i[8]
port 378 nsew signal input
rlabel metal3 s 59600 3024 59900 3080 6 wbs_dat_i[9]
port 379 nsew signal input
rlabel metal3 s 100 12096 400 12152 6 wbs_dat_o[0]
port 380 nsew signal output
rlabel metal3 s 59600 34272 59900 34328 6 wbs_dat_o[10]
port 381 nsew signal output
rlabel metal2 s 1008 100 1064 400 6 wbs_dat_o[11]
port 382 nsew signal output
rlabel metal3 s 59600 55104 59900 55160 6 wbs_dat_o[12]
port 383 nsew signal output
rlabel metal2 s 45360 59600 45416 59900 6 wbs_dat_o[13]
port 384 nsew signal output
rlabel metal3 s 59600 7056 59900 7112 6 wbs_dat_o[14]
port 385 nsew signal output
rlabel metal2 s 43008 59600 43064 59900 6 wbs_dat_o[15]
port 386 nsew signal output
rlabel metal3 s 100 16800 400 16856 6 wbs_dat_o[16]
port 387 nsew signal output
rlabel metal3 s 100 18816 400 18872 6 wbs_dat_o[17]
port 388 nsew signal output
rlabel metal2 s 40320 100 40376 400 6 wbs_dat_o[18]
port 389 nsew signal output
rlabel metal2 s 0 100 56 400 6 wbs_dat_o[19]
port 390 nsew signal output
rlabel metal2 s 47376 100 47432 400 6 wbs_dat_o[1]
port 391 nsew signal output
rlabel metal3 s 100 28224 400 28280 6 wbs_dat_o[20]
port 392 nsew signal output
rlabel metal3 s 100 52080 400 52136 6 wbs_dat_o[21]
port 393 nsew signal output
rlabel metal2 s 16128 59600 16184 59900 6 wbs_dat_o[22]
port 394 nsew signal output
rlabel metal3 s 100 19488 400 19544 6 wbs_dat_o[23]
port 395 nsew signal output
rlabel metal2 s 12432 100 12488 400 6 wbs_dat_o[24]
port 396 nsew signal output
rlabel metal2 s 4368 100 4424 400 6 wbs_dat_o[25]
port 397 nsew signal output
rlabel metal2 s 31248 59600 31304 59900 6 wbs_dat_o[26]
port 398 nsew signal output
rlabel metal2 s 17472 59600 17528 59900 6 wbs_dat_o[27]
port 399 nsew signal output
rlabel metal2 s 32256 100 32312 400 6 wbs_dat_o[28]
port 400 nsew signal output
rlabel metal2 s 41664 59600 41720 59900 6 wbs_dat_o[29]
port 401 nsew signal output
rlabel metal3 s 59600 16800 59900 16856 6 wbs_dat_o[2]
port 402 nsew signal output
rlabel metal3 s 100 39312 400 39368 6 wbs_dat_o[30]
port 403 nsew signal output
rlabel metal3 s 59600 46368 59900 46424 6 wbs_dat_o[31]
port 404 nsew signal output
rlabel metal2 s 13104 100 13160 400 6 wbs_dat_o[3]
port 405 nsew signal output
rlabel metal2 s 23184 100 23240 400 6 wbs_dat_o[4]
port 406 nsew signal output
rlabel metal3 s 100 5040 400 5096 6 wbs_dat_o[5]
port 407 nsew signal output
rlabel metal3 s 59600 44688 59900 44744 6 wbs_dat_o[6]
port 408 nsew signal output
rlabel metal2 s 36288 100 36344 400 6 wbs_dat_o[7]
port 409 nsew signal output
rlabel metal2 s 39312 59600 39368 59900 6 wbs_dat_o[8]
port 410 nsew signal output
rlabel metal2 s 38976 59600 39032 59900 6 wbs_dat_o[9]
port 411 nsew signal output
rlabel metal3 s 100 55440 400 55496 6 wbs_sel_i[0]
port 412 nsew signal input
rlabel metal2 s 6384 59600 6440 59900 6 wbs_sel_i[1]
port 413 nsew signal input
rlabel metal2 s 43344 100 43400 400 6 wbs_sel_i[2]
port 414 nsew signal input
rlabel metal3 s 100 13104 400 13160 6 wbs_sel_i[3]
port 415 nsew signal input
rlabel metal3 s 100 49728 400 49784 6 wbs_stb_i
port 416 nsew signal input
rlabel metal3 s 59600 29568 59900 29624 6 wbs_we_i
port 417 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 60000 60000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 7063522
string GDS_FILE /home/videogamo/Work/gfmpw-0/caravel_user_project/openlane/caravel_hack_soc/runs/22_12_05_18_25/results/signoff/caravel_hack_soc.magic.gds
string GDS_START 455610
<< end >>

