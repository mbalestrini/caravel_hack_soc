magic
tech gf180mcuC
magscale 1 5
timestamp 1670290645
<< obsm1 >>
rect 672 855 99288 98422
<< metal2 >>
rect 0 99600 56 99900
rect 1008 99600 1064 99900
rect 2016 99600 2072 99900
rect 3024 99600 3080 99900
rect 4032 99600 4088 99900
rect 5040 99600 5096 99900
rect 5712 99600 5768 99900
rect 6720 99600 6776 99900
rect 7728 99600 7784 99900
rect 8736 99600 8792 99900
rect 9744 99600 9800 99900
rect 10752 99600 10808 99900
rect 11760 99600 11816 99900
rect 12768 99600 12824 99900
rect 13440 99600 13496 99900
rect 14448 99600 14504 99900
rect 15456 99600 15512 99900
rect 16464 99600 16520 99900
rect 17472 99600 17528 99900
rect 18480 99600 18536 99900
rect 19488 99600 19544 99900
rect 20496 99600 20552 99900
rect 21168 99600 21224 99900
rect 22176 99600 22232 99900
rect 23184 99600 23240 99900
rect 24192 99600 24248 99900
rect 25200 99600 25256 99900
rect 26208 99600 26264 99900
rect 27216 99600 27272 99900
rect 28224 99600 28280 99900
rect 28896 99600 28952 99900
rect 29904 99600 29960 99900
rect 30912 99600 30968 99900
rect 31920 99600 31976 99900
rect 32928 99600 32984 99900
rect 33936 99600 33992 99900
rect 34944 99600 35000 99900
rect 35616 99600 35672 99900
rect 36624 99600 36680 99900
rect 37632 99600 37688 99900
rect 38640 99600 38696 99900
rect 39648 99600 39704 99900
rect 40656 99600 40712 99900
rect 41664 99600 41720 99900
rect 42672 99600 42728 99900
rect 43344 99600 43400 99900
rect 44352 99600 44408 99900
rect 45360 99600 45416 99900
rect 46368 99600 46424 99900
rect 47376 99600 47432 99900
rect 48384 99600 48440 99900
rect 49392 99600 49448 99900
rect 50400 99600 50456 99900
rect 51072 99600 51128 99900
rect 52080 99600 52136 99900
rect 53088 99600 53144 99900
rect 54096 99600 54152 99900
rect 55104 99600 55160 99900
rect 56112 99600 56168 99900
rect 57120 99600 57176 99900
rect 58128 99600 58184 99900
rect 58800 99600 58856 99900
rect 59808 99600 59864 99900
rect 60816 99600 60872 99900
rect 61824 99600 61880 99900
rect 62832 99600 62888 99900
rect 63840 99600 63896 99900
rect 64848 99600 64904 99900
rect 65856 99600 65912 99900
rect 66528 99600 66584 99900
rect 67536 99600 67592 99900
rect 68544 99600 68600 99900
rect 69552 99600 69608 99900
rect 70560 99600 70616 99900
rect 71568 99600 71624 99900
rect 72576 99600 72632 99900
rect 73584 99600 73640 99900
rect 74256 99600 74312 99900
rect 75264 99600 75320 99900
rect 76272 99600 76328 99900
rect 77280 99600 77336 99900
rect 78288 99600 78344 99900
rect 79296 99600 79352 99900
rect 80304 99600 80360 99900
rect 80976 99600 81032 99900
rect 81984 99600 82040 99900
rect 82992 99600 83048 99900
rect 84000 99600 84056 99900
rect 85008 99600 85064 99900
rect 86016 99600 86072 99900
rect 87024 99600 87080 99900
rect 88032 99600 88088 99900
rect 88704 99600 88760 99900
rect 89712 99600 89768 99900
rect 90720 99600 90776 99900
rect 91728 99600 91784 99900
rect 92736 99600 92792 99900
rect 93744 99600 93800 99900
rect 94752 99600 94808 99900
rect 95760 99600 95816 99900
rect 96432 99600 96488 99900
rect 97440 99600 97496 99900
rect 98448 99600 98504 99900
rect 99456 99600 99512 99900
rect 0 100 56 400
rect 672 100 728 400
rect 1680 100 1736 400
rect 2688 100 2744 400
rect 3696 100 3752 400
rect 4704 100 4760 400
rect 5712 100 5768 400
rect 6720 100 6776 400
rect 7392 100 7448 400
rect 8400 100 8456 400
rect 9408 100 9464 400
rect 10416 100 10472 400
rect 11424 100 11480 400
rect 12432 100 12488 400
rect 13440 100 13496 400
rect 14448 100 14504 400
rect 15120 100 15176 400
rect 16128 100 16184 400
rect 17136 100 17192 400
rect 18144 100 18200 400
rect 19152 100 19208 400
rect 20160 100 20216 400
rect 21168 100 21224 400
rect 22176 100 22232 400
rect 22848 100 22904 400
rect 23856 100 23912 400
rect 24864 100 24920 400
rect 25872 100 25928 400
rect 26880 100 26936 400
rect 27888 100 27944 400
rect 28896 100 28952 400
rect 29904 100 29960 400
rect 30576 100 30632 400
rect 31584 100 31640 400
rect 32592 100 32648 400
rect 33600 100 33656 400
rect 34608 100 34664 400
rect 35616 100 35672 400
rect 36624 100 36680 400
rect 37632 100 37688 400
rect 38304 100 38360 400
rect 39312 100 39368 400
rect 40320 100 40376 400
rect 41328 100 41384 400
rect 42336 100 42392 400
rect 43344 100 43400 400
rect 44352 100 44408 400
rect 45024 100 45080 400
rect 46032 100 46088 400
rect 47040 100 47096 400
rect 48048 100 48104 400
rect 49056 100 49112 400
rect 50064 100 50120 400
rect 51072 100 51128 400
rect 52080 100 52136 400
rect 52752 100 52808 400
rect 53760 100 53816 400
rect 54768 100 54824 400
rect 55776 100 55832 400
rect 56784 100 56840 400
rect 57792 100 57848 400
rect 58800 100 58856 400
rect 59808 100 59864 400
rect 60480 100 60536 400
rect 61488 100 61544 400
rect 62496 100 62552 400
rect 63504 100 63560 400
rect 64512 100 64568 400
rect 65520 100 65576 400
rect 66528 100 66584 400
rect 67536 100 67592 400
rect 68208 100 68264 400
rect 69216 100 69272 400
rect 70224 100 70280 400
rect 71232 100 71288 400
rect 72240 100 72296 400
rect 73248 100 73304 400
rect 74256 100 74312 400
rect 75264 100 75320 400
rect 75936 100 75992 400
rect 76944 100 77000 400
rect 77952 100 78008 400
rect 78960 100 79016 400
rect 79968 100 80024 400
rect 80976 100 81032 400
rect 81984 100 82040 400
rect 82992 100 83048 400
rect 83664 100 83720 400
rect 84672 100 84728 400
rect 85680 100 85736 400
rect 86688 100 86744 400
rect 87696 100 87752 400
rect 88704 100 88760 400
rect 89712 100 89768 400
rect 90384 100 90440 400
rect 91392 100 91448 400
rect 92400 100 92456 400
rect 93408 100 93464 400
rect 94416 100 94472 400
rect 95424 100 95480 400
rect 96432 100 96488 400
rect 97440 100 97496 400
rect 98112 100 98168 400
rect 99120 100 99176 400
<< obsm2 >>
rect 86 99570 978 99666
rect 1094 99570 1986 99666
rect 2102 99570 2994 99666
rect 3110 99570 4002 99666
rect 4118 99570 5010 99666
rect 5126 99570 5682 99666
rect 5798 99570 6690 99666
rect 6806 99570 7698 99666
rect 7814 99570 8706 99666
rect 8822 99570 9714 99666
rect 9830 99570 10722 99666
rect 10838 99570 11730 99666
rect 11846 99570 12738 99666
rect 12854 99570 13410 99666
rect 13526 99570 14418 99666
rect 14534 99570 15426 99666
rect 15542 99570 16434 99666
rect 16550 99570 17442 99666
rect 17558 99570 18450 99666
rect 18566 99570 19458 99666
rect 19574 99570 20466 99666
rect 20582 99570 21138 99666
rect 21254 99570 22146 99666
rect 22262 99570 23154 99666
rect 23270 99570 24162 99666
rect 24278 99570 25170 99666
rect 25286 99570 26178 99666
rect 26294 99570 27186 99666
rect 27302 99570 28194 99666
rect 28310 99570 28866 99666
rect 28982 99570 29874 99666
rect 29990 99570 30882 99666
rect 30998 99570 31890 99666
rect 32006 99570 32898 99666
rect 33014 99570 33906 99666
rect 34022 99570 34914 99666
rect 35030 99570 35586 99666
rect 35702 99570 36594 99666
rect 36710 99570 37602 99666
rect 37718 99570 38610 99666
rect 38726 99570 39618 99666
rect 39734 99570 40626 99666
rect 40742 99570 41634 99666
rect 41750 99570 42642 99666
rect 42758 99570 43314 99666
rect 43430 99570 44322 99666
rect 44438 99570 45330 99666
rect 45446 99570 46338 99666
rect 46454 99570 47346 99666
rect 47462 99570 48354 99666
rect 48470 99570 49362 99666
rect 49478 99570 50370 99666
rect 50486 99570 51042 99666
rect 51158 99570 52050 99666
rect 52166 99570 53058 99666
rect 53174 99570 54066 99666
rect 54182 99570 55074 99666
rect 55190 99570 56082 99666
rect 56198 99570 57090 99666
rect 57206 99570 58098 99666
rect 58214 99570 58770 99666
rect 58886 99570 59778 99666
rect 59894 99570 60786 99666
rect 60902 99570 61794 99666
rect 61910 99570 62802 99666
rect 62918 99570 63810 99666
rect 63926 99570 64818 99666
rect 64934 99570 65826 99666
rect 65942 99570 66498 99666
rect 66614 99570 67506 99666
rect 67622 99570 68514 99666
rect 68630 99570 69522 99666
rect 69638 99570 70530 99666
rect 70646 99570 71538 99666
rect 71654 99570 72546 99666
rect 72662 99570 73554 99666
rect 73670 99570 74226 99666
rect 74342 99570 75234 99666
rect 75350 99570 76242 99666
rect 76358 99570 77250 99666
rect 77366 99570 78258 99666
rect 78374 99570 79266 99666
rect 79382 99570 80274 99666
rect 80390 99570 80946 99666
rect 81062 99570 81954 99666
rect 82070 99570 82962 99666
rect 83078 99570 83970 99666
rect 84086 99570 84978 99666
rect 85094 99570 85986 99666
rect 86102 99570 86994 99666
rect 87110 99570 88002 99666
rect 88118 99570 88674 99666
rect 88790 99570 89682 99666
rect 89798 99570 90690 99666
rect 90806 99570 91698 99666
rect 91814 99570 92706 99666
rect 92822 99570 93714 99666
rect 93830 99570 94722 99666
rect 94838 99570 95730 99666
rect 95846 99570 96402 99666
rect 96518 99570 97410 99666
rect 97526 99570 98418 99666
rect 98534 99570 99050 99666
rect 14 430 99050 99570
rect 86 400 642 430
rect 758 400 1650 430
rect 1766 400 2658 430
rect 2774 400 3666 430
rect 3782 400 4674 430
rect 4790 400 5682 430
rect 5798 400 6690 430
rect 6806 400 7362 430
rect 7478 400 8370 430
rect 8486 400 9378 430
rect 9494 400 10386 430
rect 10502 400 11394 430
rect 11510 400 12402 430
rect 12518 400 13410 430
rect 13526 400 14418 430
rect 14534 400 15090 430
rect 15206 400 16098 430
rect 16214 400 17106 430
rect 17222 400 18114 430
rect 18230 400 19122 430
rect 19238 400 20130 430
rect 20246 400 21138 430
rect 21254 400 22146 430
rect 22262 400 22818 430
rect 22934 400 23826 430
rect 23942 400 24834 430
rect 24950 400 25842 430
rect 25958 400 26850 430
rect 26966 400 27858 430
rect 27974 400 28866 430
rect 28982 400 29874 430
rect 29990 400 30546 430
rect 30662 400 31554 430
rect 31670 400 32562 430
rect 32678 400 33570 430
rect 33686 400 34578 430
rect 34694 400 35586 430
rect 35702 400 36594 430
rect 36710 400 37602 430
rect 37718 400 38274 430
rect 38390 400 39282 430
rect 39398 400 40290 430
rect 40406 400 41298 430
rect 41414 400 42306 430
rect 42422 400 43314 430
rect 43430 400 44322 430
rect 44438 400 44994 430
rect 45110 400 46002 430
rect 46118 400 47010 430
rect 47126 400 48018 430
rect 48134 400 49026 430
rect 49142 400 50034 430
rect 50150 400 51042 430
rect 51158 400 52050 430
rect 52166 400 52722 430
rect 52838 400 53730 430
rect 53846 400 54738 430
rect 54854 400 55746 430
rect 55862 400 56754 430
rect 56870 400 57762 430
rect 57878 400 58770 430
rect 58886 400 59778 430
rect 59894 400 60450 430
rect 60566 400 61458 430
rect 61574 400 62466 430
rect 62582 400 63474 430
rect 63590 400 64482 430
rect 64598 400 65490 430
rect 65606 400 66498 430
rect 66614 400 67506 430
rect 67622 400 68178 430
rect 68294 400 69186 430
rect 69302 400 70194 430
rect 70310 400 71202 430
rect 71318 400 72210 430
rect 72326 400 73218 430
rect 73334 400 74226 430
rect 74342 400 75234 430
rect 75350 400 75906 430
rect 76022 400 76914 430
rect 77030 400 77922 430
rect 78038 400 78930 430
rect 79046 400 79938 430
rect 80054 400 80946 430
rect 81062 400 81954 430
rect 82070 400 82962 430
rect 83078 400 83634 430
rect 83750 400 84642 430
rect 84758 400 85650 430
rect 85766 400 86658 430
rect 86774 400 87666 430
rect 87782 400 88674 430
rect 88790 400 89682 430
rect 89798 400 90354 430
rect 90470 400 91362 430
rect 91478 400 92370 430
rect 92486 400 93378 430
rect 93494 400 94386 430
rect 94502 400 95394 430
rect 95510 400 96402 430
rect 96518 400 97410 430
rect 97526 400 98082 430
rect 98198 400 99050 430
<< metal3 >>
rect 99600 99456 99900 99512
rect 100 99120 400 99176
rect 99600 98448 99900 98504
rect 100 98112 400 98168
rect 100 97440 400 97496
rect 99600 97440 99900 97496
rect 100 96432 400 96488
rect 99600 96432 99900 96488
rect 99600 95760 99900 95816
rect 100 95424 400 95480
rect 99600 94752 99900 94808
rect 100 94416 400 94472
rect 99600 93744 99900 93800
rect 100 93408 400 93464
rect 99600 92736 99900 92792
rect 100 92400 400 92456
rect 99600 91728 99900 91784
rect 100 91392 400 91448
rect 99600 90720 99900 90776
rect 100 90384 400 90440
rect 100 89712 400 89768
rect 99600 89712 99900 89768
rect 100 88704 400 88760
rect 99600 88704 99900 88760
rect 99600 88032 99900 88088
rect 100 87696 400 87752
rect 99600 87024 99900 87080
rect 100 86688 400 86744
rect 99600 86016 99900 86072
rect 100 85680 400 85736
rect 99600 85008 99900 85064
rect 100 84672 400 84728
rect 99600 84000 99900 84056
rect 100 83664 400 83720
rect 100 82992 400 83048
rect 99600 82992 99900 83048
rect 100 81984 400 82040
rect 99600 81984 99900 82040
rect 100 80976 400 81032
rect 99600 80976 99900 81032
rect 99600 80304 99900 80360
rect 100 79968 400 80024
rect 99600 79296 99900 79352
rect 100 78960 400 79016
rect 99600 78288 99900 78344
rect 100 77952 400 78008
rect 99600 77280 99900 77336
rect 100 76944 400 77000
rect 99600 76272 99900 76328
rect 100 75936 400 75992
rect 100 75264 400 75320
rect 99600 75264 99900 75320
rect 100 74256 400 74312
rect 99600 74256 99900 74312
rect 99600 73584 99900 73640
rect 100 73248 400 73304
rect 99600 72576 99900 72632
rect 100 72240 400 72296
rect 99600 71568 99900 71624
rect 100 71232 400 71288
rect 99600 70560 99900 70616
rect 100 70224 400 70280
rect 99600 69552 99900 69608
rect 100 69216 400 69272
rect 99600 68544 99900 68600
rect 100 68208 400 68264
rect 100 67536 400 67592
rect 99600 67536 99900 67592
rect 100 66528 400 66584
rect 99600 66528 99900 66584
rect 99600 65856 99900 65912
rect 100 65520 400 65576
rect 99600 64848 99900 64904
rect 100 64512 400 64568
rect 99600 63840 99900 63896
rect 100 63504 400 63560
rect 99600 62832 99900 62888
rect 100 62496 400 62552
rect 99600 61824 99900 61880
rect 100 61488 400 61544
rect 99600 60816 99900 60872
rect 100 60480 400 60536
rect 100 59808 400 59864
rect 99600 59808 99900 59864
rect 100 58800 400 58856
rect 99600 58800 99900 58856
rect 99600 58128 99900 58184
rect 100 57792 400 57848
rect 99600 57120 99900 57176
rect 100 56784 400 56840
rect 99600 56112 99900 56168
rect 100 55776 400 55832
rect 99600 55104 99900 55160
rect 100 54768 400 54824
rect 99600 54096 99900 54152
rect 100 53760 400 53816
rect 99600 53088 99900 53144
rect 100 52752 400 52808
rect 100 52080 400 52136
rect 99600 52080 99900 52136
rect 100 51072 400 51128
rect 99600 51072 99900 51128
rect 99600 50400 99900 50456
rect 100 50064 400 50120
rect 99600 49392 99900 49448
rect 100 49056 400 49112
rect 99600 48384 99900 48440
rect 100 48048 400 48104
rect 99600 47376 99900 47432
rect 100 47040 400 47096
rect 99600 46368 99900 46424
rect 100 46032 400 46088
rect 99600 45360 99900 45416
rect 100 45024 400 45080
rect 100 44352 400 44408
rect 99600 44352 99900 44408
rect 100 43344 400 43400
rect 99600 43344 99900 43400
rect 99600 42672 99900 42728
rect 100 42336 400 42392
rect 99600 41664 99900 41720
rect 100 41328 400 41384
rect 99600 40656 99900 40712
rect 100 40320 400 40376
rect 99600 39648 99900 39704
rect 100 39312 400 39368
rect 99600 38640 99900 38696
rect 100 38304 400 38360
rect 100 37632 400 37688
rect 99600 37632 99900 37688
rect 100 36624 400 36680
rect 99600 36624 99900 36680
rect 100 35616 400 35672
rect 99600 35616 99900 35672
rect 99600 34944 99900 35000
rect 100 34608 400 34664
rect 99600 33936 99900 33992
rect 100 33600 400 33656
rect 99600 32928 99900 32984
rect 100 32592 400 32648
rect 99600 31920 99900 31976
rect 100 31584 400 31640
rect 99600 30912 99900 30968
rect 100 30576 400 30632
rect 100 29904 400 29960
rect 99600 29904 99900 29960
rect 100 28896 400 28952
rect 99600 28896 99900 28952
rect 99600 28224 99900 28280
rect 100 27888 400 27944
rect 99600 27216 99900 27272
rect 100 26880 400 26936
rect 99600 26208 99900 26264
rect 100 25872 400 25928
rect 99600 25200 99900 25256
rect 100 24864 400 24920
rect 99600 24192 99900 24248
rect 100 23856 400 23912
rect 99600 23184 99900 23240
rect 100 22848 400 22904
rect 100 22176 400 22232
rect 99600 22176 99900 22232
rect 100 21168 400 21224
rect 99600 21168 99900 21224
rect 99600 20496 99900 20552
rect 100 20160 400 20216
rect 99600 19488 99900 19544
rect 100 19152 400 19208
rect 99600 18480 99900 18536
rect 100 18144 400 18200
rect 99600 17472 99900 17528
rect 100 17136 400 17192
rect 99600 16464 99900 16520
rect 100 16128 400 16184
rect 99600 15456 99900 15512
rect 100 15120 400 15176
rect 100 14448 400 14504
rect 99600 14448 99900 14504
rect 100 13440 400 13496
rect 99600 13440 99900 13496
rect 99600 12768 99900 12824
rect 100 12432 400 12488
rect 99600 11760 99900 11816
rect 100 11424 400 11480
rect 99600 10752 99900 10808
rect 100 10416 400 10472
rect 99600 9744 99900 9800
rect 100 9408 400 9464
rect 99600 8736 99900 8792
rect 100 8400 400 8456
rect 99600 7728 99900 7784
rect 100 7392 400 7448
rect 100 6720 400 6776
rect 99600 6720 99900 6776
rect 100 5712 400 5768
rect 99600 5712 99900 5768
rect 99600 5040 99900 5096
rect 100 4704 400 4760
rect 99600 4032 99900 4088
rect 100 3696 400 3752
rect 99600 3024 99900 3080
rect 100 2688 400 2744
rect 99600 2016 99900 2072
rect 100 1680 400 1736
rect 99600 1008 99900 1064
rect 100 672 400 728
rect 99600 0 99900 56
<< obsm3 >>
rect 9 99426 99570 99498
rect 9 99206 99666 99426
rect 9 99090 70 99206
rect 430 99090 99666 99206
rect 9 98534 99666 99090
rect 9 98418 99570 98534
rect 9 98198 99666 98418
rect 9 98082 70 98198
rect 430 98082 99666 98198
rect 9 97526 99666 98082
rect 9 97410 70 97526
rect 430 97410 99570 97526
rect 9 96518 99666 97410
rect 9 96402 70 96518
rect 430 96402 99570 96518
rect 9 95846 99666 96402
rect 9 95730 99570 95846
rect 9 95510 99666 95730
rect 9 95394 70 95510
rect 430 95394 99666 95510
rect 9 94838 99666 95394
rect 9 94722 99570 94838
rect 9 94502 99666 94722
rect 9 94386 70 94502
rect 430 94386 99666 94502
rect 9 93830 99666 94386
rect 9 93714 99570 93830
rect 9 93494 99666 93714
rect 9 93378 70 93494
rect 430 93378 99666 93494
rect 9 92822 99666 93378
rect 9 92706 99570 92822
rect 9 92486 99666 92706
rect 9 92370 70 92486
rect 430 92370 99666 92486
rect 9 91814 99666 92370
rect 9 91698 99570 91814
rect 9 91478 99666 91698
rect 9 91362 70 91478
rect 430 91362 99666 91478
rect 9 90806 99666 91362
rect 9 90690 99570 90806
rect 9 90470 99666 90690
rect 9 90354 70 90470
rect 430 90354 99666 90470
rect 9 89798 99666 90354
rect 9 89682 70 89798
rect 430 89682 99570 89798
rect 9 88790 99666 89682
rect 9 88674 70 88790
rect 430 88674 99570 88790
rect 9 88118 99666 88674
rect 9 88002 99570 88118
rect 9 87782 99666 88002
rect 9 87666 70 87782
rect 430 87666 99666 87782
rect 9 87110 99666 87666
rect 9 86994 99570 87110
rect 9 86774 99666 86994
rect 9 86658 70 86774
rect 430 86658 99666 86774
rect 9 86102 99666 86658
rect 9 85986 99570 86102
rect 9 85766 99666 85986
rect 9 85650 70 85766
rect 430 85650 99666 85766
rect 9 85094 99666 85650
rect 9 84978 99570 85094
rect 9 84758 99666 84978
rect 9 84642 70 84758
rect 430 84642 99666 84758
rect 9 84086 99666 84642
rect 9 83970 99570 84086
rect 9 83750 99666 83970
rect 9 83634 70 83750
rect 430 83634 99666 83750
rect 9 83078 99666 83634
rect 9 82962 70 83078
rect 430 82962 99570 83078
rect 9 82070 99666 82962
rect 9 81954 70 82070
rect 430 81954 99570 82070
rect 9 81062 99666 81954
rect 9 80946 70 81062
rect 430 80946 99570 81062
rect 9 80390 99666 80946
rect 9 80274 99570 80390
rect 9 80054 99666 80274
rect 9 79938 70 80054
rect 430 79938 99666 80054
rect 9 79382 99666 79938
rect 9 79266 99570 79382
rect 9 79046 99666 79266
rect 9 78930 70 79046
rect 430 78930 99666 79046
rect 9 78374 99666 78930
rect 9 78258 99570 78374
rect 9 78038 99666 78258
rect 9 77922 70 78038
rect 430 77922 99666 78038
rect 9 77366 99666 77922
rect 9 77250 99570 77366
rect 9 77030 99666 77250
rect 9 76914 70 77030
rect 430 76914 99666 77030
rect 9 76358 99666 76914
rect 9 76242 99570 76358
rect 9 76022 99666 76242
rect 9 75906 70 76022
rect 430 75906 99666 76022
rect 9 75350 99666 75906
rect 9 75234 70 75350
rect 430 75234 99570 75350
rect 9 74342 99666 75234
rect 9 74226 70 74342
rect 430 74226 99570 74342
rect 9 73670 99666 74226
rect 9 73554 99570 73670
rect 9 73334 99666 73554
rect 9 73218 70 73334
rect 430 73218 99666 73334
rect 9 72662 99666 73218
rect 9 72546 99570 72662
rect 9 72326 99666 72546
rect 9 72210 70 72326
rect 430 72210 99666 72326
rect 9 71654 99666 72210
rect 9 71538 99570 71654
rect 9 71318 99666 71538
rect 9 71202 70 71318
rect 430 71202 99666 71318
rect 9 70646 99666 71202
rect 9 70530 99570 70646
rect 9 70310 99666 70530
rect 9 70194 70 70310
rect 430 70194 99666 70310
rect 9 69638 99666 70194
rect 9 69522 99570 69638
rect 9 69302 99666 69522
rect 9 69186 70 69302
rect 430 69186 99666 69302
rect 9 68630 99666 69186
rect 9 68514 99570 68630
rect 9 68294 99666 68514
rect 9 68178 70 68294
rect 430 68178 99666 68294
rect 9 67622 99666 68178
rect 9 67506 70 67622
rect 430 67506 99570 67622
rect 9 66614 99666 67506
rect 9 66498 70 66614
rect 430 66498 99570 66614
rect 9 65942 99666 66498
rect 9 65826 99570 65942
rect 9 65606 99666 65826
rect 9 65490 70 65606
rect 430 65490 99666 65606
rect 9 64934 99666 65490
rect 9 64818 99570 64934
rect 9 64598 99666 64818
rect 9 64482 70 64598
rect 430 64482 99666 64598
rect 9 63926 99666 64482
rect 9 63810 99570 63926
rect 9 63590 99666 63810
rect 9 63474 70 63590
rect 430 63474 99666 63590
rect 9 62918 99666 63474
rect 9 62802 99570 62918
rect 9 62582 99666 62802
rect 9 62466 70 62582
rect 430 62466 99666 62582
rect 9 61910 99666 62466
rect 9 61794 99570 61910
rect 9 61574 99666 61794
rect 9 61458 70 61574
rect 430 61458 99666 61574
rect 9 60902 99666 61458
rect 9 60786 99570 60902
rect 9 60566 99666 60786
rect 9 60450 70 60566
rect 430 60450 99666 60566
rect 9 59894 99666 60450
rect 9 59778 70 59894
rect 430 59778 99570 59894
rect 9 58886 99666 59778
rect 9 58770 70 58886
rect 430 58770 99570 58886
rect 9 58214 99666 58770
rect 9 58098 99570 58214
rect 9 57878 99666 58098
rect 9 57762 70 57878
rect 430 57762 99666 57878
rect 9 57206 99666 57762
rect 9 57090 99570 57206
rect 9 56870 99666 57090
rect 9 56754 70 56870
rect 430 56754 99666 56870
rect 9 56198 99666 56754
rect 9 56082 99570 56198
rect 9 55862 99666 56082
rect 9 55746 70 55862
rect 430 55746 99666 55862
rect 9 55190 99666 55746
rect 9 55074 99570 55190
rect 9 54854 99666 55074
rect 9 54738 70 54854
rect 430 54738 99666 54854
rect 9 54182 99666 54738
rect 9 54066 99570 54182
rect 9 53846 99666 54066
rect 9 53730 70 53846
rect 430 53730 99666 53846
rect 9 53174 99666 53730
rect 9 53058 99570 53174
rect 9 52838 99666 53058
rect 9 52722 70 52838
rect 430 52722 99666 52838
rect 9 52166 99666 52722
rect 9 52050 70 52166
rect 430 52050 99570 52166
rect 9 51158 99666 52050
rect 9 51042 70 51158
rect 430 51042 99570 51158
rect 9 50486 99666 51042
rect 9 50370 99570 50486
rect 9 50150 99666 50370
rect 9 50034 70 50150
rect 430 50034 99666 50150
rect 9 49478 99666 50034
rect 9 49362 99570 49478
rect 9 49142 99666 49362
rect 9 49026 70 49142
rect 430 49026 99666 49142
rect 9 48470 99666 49026
rect 9 48354 99570 48470
rect 9 48134 99666 48354
rect 9 48018 70 48134
rect 430 48018 99666 48134
rect 9 47462 99666 48018
rect 9 47346 99570 47462
rect 9 47126 99666 47346
rect 9 47010 70 47126
rect 430 47010 99666 47126
rect 9 46454 99666 47010
rect 9 46338 99570 46454
rect 9 46118 99666 46338
rect 9 46002 70 46118
rect 430 46002 99666 46118
rect 9 45446 99666 46002
rect 9 45330 99570 45446
rect 9 45110 99666 45330
rect 9 44994 70 45110
rect 430 44994 99666 45110
rect 9 44438 99666 44994
rect 9 44322 70 44438
rect 430 44322 99570 44438
rect 9 43430 99666 44322
rect 9 43314 70 43430
rect 430 43314 99570 43430
rect 9 42758 99666 43314
rect 9 42642 99570 42758
rect 9 42422 99666 42642
rect 9 42306 70 42422
rect 430 42306 99666 42422
rect 9 41750 99666 42306
rect 9 41634 99570 41750
rect 9 41414 99666 41634
rect 9 41298 70 41414
rect 430 41298 99666 41414
rect 9 40742 99666 41298
rect 9 40626 99570 40742
rect 9 40406 99666 40626
rect 9 40290 70 40406
rect 430 40290 99666 40406
rect 9 39734 99666 40290
rect 9 39618 99570 39734
rect 9 39398 99666 39618
rect 9 39282 70 39398
rect 430 39282 99666 39398
rect 9 38726 99666 39282
rect 9 38610 99570 38726
rect 9 38390 99666 38610
rect 9 38274 70 38390
rect 430 38274 99666 38390
rect 9 37718 99666 38274
rect 9 37602 70 37718
rect 430 37602 99570 37718
rect 9 36710 99666 37602
rect 9 36594 70 36710
rect 430 36594 99570 36710
rect 9 35702 99666 36594
rect 9 35586 70 35702
rect 430 35586 99570 35702
rect 9 35030 99666 35586
rect 9 34914 99570 35030
rect 9 34694 99666 34914
rect 9 34578 70 34694
rect 430 34578 99666 34694
rect 9 34022 99666 34578
rect 9 33906 99570 34022
rect 9 33686 99666 33906
rect 9 33570 70 33686
rect 430 33570 99666 33686
rect 9 33014 99666 33570
rect 9 32898 99570 33014
rect 9 32678 99666 32898
rect 9 32562 70 32678
rect 430 32562 99666 32678
rect 9 32006 99666 32562
rect 9 31890 99570 32006
rect 9 31670 99666 31890
rect 9 31554 70 31670
rect 430 31554 99666 31670
rect 9 30998 99666 31554
rect 9 30882 99570 30998
rect 9 30662 99666 30882
rect 9 30546 70 30662
rect 430 30546 99666 30662
rect 9 29990 99666 30546
rect 9 29874 70 29990
rect 430 29874 99570 29990
rect 9 28982 99666 29874
rect 9 28866 70 28982
rect 430 28866 99570 28982
rect 9 28310 99666 28866
rect 9 28194 99570 28310
rect 9 27974 99666 28194
rect 9 27858 70 27974
rect 430 27858 99666 27974
rect 9 27302 99666 27858
rect 9 27186 99570 27302
rect 9 26966 99666 27186
rect 9 26850 70 26966
rect 430 26850 99666 26966
rect 9 26294 99666 26850
rect 9 26178 99570 26294
rect 9 25958 99666 26178
rect 9 25842 70 25958
rect 430 25842 99666 25958
rect 9 25286 99666 25842
rect 9 25170 99570 25286
rect 9 24950 99666 25170
rect 9 24834 70 24950
rect 430 24834 99666 24950
rect 9 24278 99666 24834
rect 9 24162 99570 24278
rect 9 23942 99666 24162
rect 9 23826 70 23942
rect 430 23826 99666 23942
rect 9 23270 99666 23826
rect 9 23154 99570 23270
rect 9 22934 99666 23154
rect 9 22818 70 22934
rect 430 22818 99666 22934
rect 9 22262 99666 22818
rect 9 22146 70 22262
rect 430 22146 99570 22262
rect 9 21254 99666 22146
rect 9 21138 70 21254
rect 430 21138 99570 21254
rect 9 20582 99666 21138
rect 9 20466 99570 20582
rect 9 20246 99666 20466
rect 9 20130 70 20246
rect 430 20130 99666 20246
rect 9 19574 99666 20130
rect 9 19458 99570 19574
rect 9 19238 99666 19458
rect 9 19122 70 19238
rect 430 19122 99666 19238
rect 9 18566 99666 19122
rect 9 18450 99570 18566
rect 9 18230 99666 18450
rect 9 18114 70 18230
rect 430 18114 99666 18230
rect 9 17558 99666 18114
rect 9 17442 99570 17558
rect 9 17222 99666 17442
rect 9 17106 70 17222
rect 430 17106 99666 17222
rect 9 16550 99666 17106
rect 9 16434 99570 16550
rect 9 16214 99666 16434
rect 9 16098 70 16214
rect 430 16098 99666 16214
rect 9 15542 99666 16098
rect 9 15426 99570 15542
rect 9 15206 99666 15426
rect 9 15090 70 15206
rect 430 15090 99666 15206
rect 9 14534 99666 15090
rect 9 14418 70 14534
rect 430 14418 99570 14534
rect 9 13526 99666 14418
rect 9 13410 70 13526
rect 430 13410 99570 13526
rect 9 12854 99666 13410
rect 9 12738 99570 12854
rect 9 12518 99666 12738
rect 9 12402 70 12518
rect 430 12402 99666 12518
rect 9 11846 99666 12402
rect 9 11730 99570 11846
rect 9 11510 99666 11730
rect 9 11394 70 11510
rect 430 11394 99666 11510
rect 9 10838 99666 11394
rect 9 10722 99570 10838
rect 9 10502 99666 10722
rect 9 10386 70 10502
rect 430 10386 99666 10502
rect 9 9830 99666 10386
rect 9 9714 99570 9830
rect 9 9494 99666 9714
rect 9 9378 70 9494
rect 430 9378 99666 9494
rect 9 8822 99666 9378
rect 9 8706 99570 8822
rect 9 8486 99666 8706
rect 9 8370 70 8486
rect 430 8370 99666 8486
rect 9 7814 99666 8370
rect 9 7698 99570 7814
rect 9 7478 99666 7698
rect 9 7362 70 7478
rect 430 7362 99666 7478
rect 9 6806 99666 7362
rect 9 6690 70 6806
rect 430 6690 99570 6806
rect 9 5798 99666 6690
rect 9 5682 70 5798
rect 430 5682 99570 5798
rect 9 5126 99666 5682
rect 9 5010 99570 5126
rect 9 4790 99666 5010
rect 9 4674 70 4790
rect 430 4674 99666 4790
rect 9 4118 99666 4674
rect 9 4002 99570 4118
rect 9 3782 99666 4002
rect 9 3666 70 3782
rect 430 3666 99666 3782
rect 9 3110 99666 3666
rect 9 2994 99570 3110
rect 9 2774 99666 2994
rect 9 2658 70 2774
rect 430 2658 99666 2774
rect 9 2102 99666 2658
rect 9 1986 99570 2102
rect 9 1766 99666 1986
rect 9 1650 70 1766
rect 430 1650 99666 1766
rect 9 1094 99666 1650
rect 9 978 99570 1094
rect 9 758 99666 978
rect 9 686 70 758
rect 430 686 99666 758
<< metal4 >>
rect 2224 1538 2384 98422
rect 9904 1538 10064 98422
rect 17584 1538 17744 98422
rect 25264 1538 25424 98422
rect 32944 1538 33104 98422
rect 40624 1538 40784 98422
rect 48304 1538 48464 98422
rect 55984 1538 56144 98422
rect 63664 1538 63824 98422
rect 71344 1538 71504 98422
rect 79024 1538 79184 98422
rect 86704 1538 86864 98422
rect 94384 1538 94544 98422
<< obsm4 >>
rect 1190 1745 2194 98271
rect 2414 1745 9874 98271
rect 10094 1745 17554 98271
rect 17774 1745 25234 98271
rect 25454 1745 32914 98271
rect 33134 1745 40594 98271
rect 40814 1745 48274 98271
rect 48494 1745 55954 98271
rect 56174 1745 63634 98271
rect 63854 1745 71314 98271
rect 71534 1745 78994 98271
rect 79214 1745 86674 98271
rect 86894 1745 87066 98271
<< obsm5 >>
rect 1182 7566 79906 69602
<< labels >>
rlabel metal3 s 100 34608 400 34664 6 io_in[0]
port 1 nsew signal input
rlabel metal3 s 100 46032 400 46088 6 io_in[10]
port 2 nsew signal input
rlabel metal3 s 100 41328 400 41384 6 io_in[11]
port 3 nsew signal input
rlabel metal2 s 96432 99600 96488 99900 6 io_in[12]
port 4 nsew signal input
rlabel metal3 s 100 35616 400 35672 6 io_in[13]
port 5 nsew signal input
rlabel metal2 s 55104 99600 55160 99900 6 io_in[14]
port 6 nsew signal input
rlabel metal3 s 99600 19488 99900 19544 6 io_in[15]
port 7 nsew signal input
rlabel metal2 s 28896 100 28952 400 6 io_in[16]
port 8 nsew signal input
rlabel metal2 s 22176 99600 22232 99900 6 io_in[17]
port 9 nsew signal input
rlabel metal3 s 100 44352 400 44408 6 io_in[18]
port 10 nsew signal input
rlabel metal3 s 99600 99456 99900 99512 6 io_in[19]
port 11 nsew signal input
rlabel metal2 s 80304 99600 80360 99900 6 io_in[1]
port 12 nsew signal input
rlabel metal2 s 58128 99600 58184 99900 6 io_in[20]
port 13 nsew signal input
rlabel metal2 s 94752 99600 94808 99900 6 io_in[21]
port 14 nsew signal input
rlabel metal2 s 2016 99600 2072 99900 6 io_in[22]
port 15 nsew signal input
rlabel metal2 s 13440 100 13496 400 6 io_in[23]
port 16 nsew signal input
rlabel metal2 s 12768 99600 12824 99900 6 io_in[24]
port 17 nsew signal input
rlabel metal2 s 16464 99600 16520 99900 6 io_in[25]
port 18 nsew signal input
rlabel metal3 s 99600 10752 99900 10808 6 io_in[26]
port 19 nsew signal input
rlabel metal3 s 100 23856 400 23912 6 io_in[27]
port 20 nsew signal input
rlabel metal2 s 4032 99600 4088 99900 6 io_in[28]
port 21 nsew signal input
rlabel metal3 s 99600 97440 99900 97496 6 io_in[29]
port 22 nsew signal input
rlabel metal3 s 100 10416 400 10472 6 io_in[2]
port 23 nsew signal input
rlabel metal2 s 70224 100 70280 400 6 io_in[30]
port 24 nsew signal input
rlabel metal2 s 14448 99600 14504 99900 6 io_in[31]
port 25 nsew signal input
rlabel metal2 s 59808 100 59864 400 6 io_in[32]
port 26 nsew signal input
rlabel metal3 s 100 98112 400 98168 6 io_in[33]
port 27 nsew signal input
rlabel metal2 s 89712 99600 89768 99900 6 io_in[34]
port 28 nsew signal input
rlabel metal2 s 21168 99600 21224 99900 6 io_in[35]
port 29 nsew signal input
rlabel metal3 s 100 25872 400 25928 6 io_in[36]
port 30 nsew signal input
rlabel metal3 s 99600 16464 99900 16520 6 io_in[37]
port 31 nsew signal input
rlabel metal3 s 100 42336 400 42392 6 io_in[3]
port 32 nsew signal input
rlabel metal2 s 89712 100 89768 400 6 io_in[4]
port 33 nsew signal input
rlabel metal3 s 100 97440 400 97496 6 io_in[5]
port 34 nsew signal input
rlabel metal3 s 100 22848 400 22904 6 io_in[6]
port 35 nsew signal input
rlabel metal3 s 99600 26208 99900 26264 6 io_in[7]
port 36 nsew signal input
rlabel metal2 s 97440 100 97496 400 6 io_in[8]
port 37 nsew signal input
rlabel metal2 s 85008 99600 85064 99900 6 io_in[9]
port 38 nsew signal input
rlabel metal2 s 3024 99600 3080 99900 6 io_oeb[0]
port 39 nsew signal output
rlabel metal3 s 100 68208 400 68264 6 io_oeb[10]
port 40 nsew signal output
rlabel metal3 s 100 62496 400 62552 6 io_oeb[11]
port 41 nsew signal output
rlabel metal3 s 100 75264 400 75320 6 io_oeb[12]
port 42 nsew signal output
rlabel metal2 s 85680 100 85736 400 6 io_oeb[13]
port 43 nsew signal output
rlabel metal2 s 98112 100 98168 400 6 io_oeb[14]
port 44 nsew signal output
rlabel metal2 s 53088 99600 53144 99900 6 io_oeb[15]
port 45 nsew signal output
rlabel metal3 s 100 57792 400 57848 6 io_oeb[16]
port 46 nsew signal output
rlabel metal2 s 9744 99600 9800 99900 6 io_oeb[17]
port 47 nsew signal output
rlabel metal3 s 100 78960 400 79016 6 io_oeb[18]
port 48 nsew signal output
rlabel metal2 s 40320 100 40376 400 6 io_oeb[19]
port 49 nsew signal output
rlabel metal3 s 99600 7728 99900 7784 6 io_oeb[1]
port 50 nsew signal output
rlabel metal2 s 84672 100 84728 400 6 io_oeb[20]
port 51 nsew signal output
rlabel metal2 s 9408 100 9464 400 6 io_oeb[21]
port 52 nsew signal output
rlabel metal3 s 99600 25200 99900 25256 6 io_oeb[22]
port 53 nsew signal output
rlabel metal3 s 100 9408 400 9464 6 io_oeb[23]
port 54 nsew signal output
rlabel metal3 s 99600 22176 99900 22232 6 io_oeb[24]
port 55 nsew signal output
rlabel metal2 s 35616 100 35672 400 6 io_oeb[25]
port 56 nsew signal output
rlabel metal2 s 82992 100 83048 400 6 io_oeb[26]
port 57 nsew signal output
rlabel metal3 s 100 66528 400 66584 6 io_oeb[27]
port 58 nsew signal output
rlabel metal3 s 100 93408 400 93464 6 io_oeb[28]
port 59 nsew signal output
rlabel metal2 s 20496 99600 20552 99900 6 io_oeb[29]
port 60 nsew signal output
rlabel metal2 s 64512 100 64568 400 6 io_oeb[2]
port 61 nsew signal output
rlabel metal3 s 100 3696 400 3752 6 io_oeb[30]
port 62 nsew signal output
rlabel metal3 s 99600 69552 99900 69608 6 io_oeb[31]
port 63 nsew signal output
rlabel metal3 s 99600 15456 99900 15512 6 io_oeb[32]
port 64 nsew signal output
rlabel metal3 s 100 81984 400 82040 6 io_oeb[33]
port 65 nsew signal output
rlabel metal3 s 100 38304 400 38360 6 io_oeb[34]
port 66 nsew signal output
rlabel metal2 s 56112 99600 56168 99900 6 io_oeb[35]
port 67 nsew signal output
rlabel metal2 s 93408 100 93464 400 6 io_oeb[36]
port 68 nsew signal output
rlabel metal3 s 100 83664 400 83720 6 io_oeb[37]
port 69 nsew signal output
rlabel metal3 s 99600 33936 99900 33992 6 io_oeb[3]
port 70 nsew signal output
rlabel metal2 s 0 99600 56 99900 6 io_oeb[4]
port 71 nsew signal output
rlabel metal3 s 99600 96432 99900 96488 6 io_oeb[5]
port 72 nsew signal output
rlabel metal2 s 48384 99600 48440 99900 6 io_oeb[6]
port 73 nsew signal output
rlabel metal3 s 99600 5712 99900 5768 6 io_oeb[7]
port 74 nsew signal output
rlabel metal3 s 99600 40656 99900 40712 6 io_oeb[8]
port 75 nsew signal output
rlabel metal3 s 99600 39648 99900 39704 6 io_oeb[9]
port 76 nsew signal output
rlabel metal3 s 100 19152 400 19208 6 io_out[0]
port 77 nsew signal output
rlabel metal2 s 97440 99600 97496 99900 6 io_out[10]
port 78 nsew signal output
rlabel metal3 s 99600 88032 99900 88088 6 io_out[11]
port 79 nsew signal output
rlabel metal3 s 99600 98448 99900 98504 6 io_out[12]
port 80 nsew signal output
rlabel metal3 s 100 74256 400 74312 6 io_out[13]
port 81 nsew signal output
rlabel metal2 s 39312 100 39368 400 6 io_out[14]
port 82 nsew signal output
rlabel metal3 s 99600 82992 99900 83048 6 io_out[15]
port 83 nsew signal output
rlabel metal2 s 11424 100 11480 400 6 io_out[16]
port 84 nsew signal output
rlabel metal2 s 83664 100 83720 400 6 io_out[17]
port 85 nsew signal output
rlabel metal2 s 65520 100 65576 400 6 io_out[18]
port 86 nsew signal output
rlabel metal2 s 6720 100 6776 400 6 io_out[19]
port 87 nsew signal output
rlabel metal2 s 68208 100 68264 400 6 io_out[1]
port 88 nsew signal output
rlabel metal2 s 45024 100 45080 400 6 io_out[20]
port 89 nsew signal output
rlabel metal2 s 33600 100 33656 400 6 io_out[21]
port 90 nsew signal output
rlabel metal3 s 100 13440 400 13496 6 io_out[22]
port 91 nsew signal output
rlabel metal2 s 73584 99600 73640 99900 6 io_out[23]
port 92 nsew signal output
rlabel metal2 s 46368 99600 46424 99900 6 io_out[24]
port 93 nsew signal output
rlabel metal2 s 42336 100 42392 400 6 io_out[25]
port 94 nsew signal output
rlabel metal2 s 70560 99600 70616 99900 6 io_out[26]
port 95 nsew signal output
rlabel metal2 s 74256 100 74312 400 6 io_out[27]
port 96 nsew signal output
rlabel metal2 s 63840 99600 63896 99900 6 io_out[28]
port 97 nsew signal output
rlabel metal2 s 94416 100 94472 400 6 io_out[29]
port 98 nsew signal output
rlabel metal2 s 91728 99600 91784 99900 6 io_out[2]
port 99 nsew signal output
rlabel metal3 s 99600 21168 99900 21224 6 io_out[30]
port 100 nsew signal output
rlabel metal2 s 84000 99600 84056 99900 6 io_out[31]
port 101 nsew signal output
rlabel metal3 s 99600 31920 99900 31976 6 io_out[32]
port 102 nsew signal output
rlabel metal2 s 66528 100 66584 400 6 io_out[33]
port 103 nsew signal output
rlabel metal3 s 99600 64848 99900 64904 6 io_out[34]
port 104 nsew signal output
rlabel metal2 s 23856 100 23912 400 6 io_out[35]
port 105 nsew signal output
rlabel metal3 s 99600 93744 99900 93800 6 io_out[36]
port 106 nsew signal output
rlabel metal3 s 99600 92736 99900 92792 6 io_out[37]
port 107 nsew signal output
rlabel metal3 s 99600 71568 99900 71624 6 io_out[3]
port 108 nsew signal output
rlabel metal3 s 100 2688 400 2744 6 io_out[4]
port 109 nsew signal output
rlabel metal3 s 100 4704 400 4760 6 io_out[5]
port 110 nsew signal output
rlabel metal3 s 100 56784 400 56840 6 io_out[6]
port 111 nsew signal output
rlabel metal2 s 62832 99600 62888 99900 6 io_out[7]
port 112 nsew signal output
rlabel metal2 s 25872 100 25928 400 6 io_out[8]
port 113 nsew signal output
rlabel metal3 s 100 51072 400 51128 6 io_out[9]
port 114 nsew signal output
rlabel metal3 s 100 70224 400 70280 6 irq[0]
port 115 nsew signal output
rlabel metal3 s 100 40320 400 40376 6 irq[1]
port 116 nsew signal output
rlabel metal2 s 30576 100 30632 400 6 irq[2]
port 117 nsew signal output
rlabel metal2 s 40656 99600 40712 99900 6 la_data_in[0]
port 118 nsew signal input
rlabel metal2 s 93744 99600 93800 99900 6 la_data_in[10]
port 119 nsew signal input
rlabel metal2 s 47040 100 47096 400 6 la_data_in[11]
port 120 nsew signal input
rlabel metal3 s 100 60480 400 60536 6 la_data_in[12]
port 121 nsew signal input
rlabel metal3 s 99600 14448 99900 14504 6 la_data_in[13]
port 122 nsew signal input
rlabel metal3 s 99600 36624 99900 36680 6 la_data_in[14]
port 123 nsew signal input
rlabel metal3 s 100 69216 400 69272 6 la_data_in[15]
port 124 nsew signal input
rlabel metal2 s 23184 99600 23240 99900 6 la_data_in[16]
port 125 nsew signal input
rlabel metal3 s 99600 20496 99900 20552 6 la_data_in[17]
port 126 nsew signal input
rlabel metal3 s 99600 75264 99900 75320 6 la_data_in[18]
port 127 nsew signal input
rlabel metal3 s 99600 44352 99900 44408 6 la_data_in[19]
port 128 nsew signal input
rlabel metal2 s 76272 99600 76328 99900 6 la_data_in[1]
port 129 nsew signal input
rlabel metal2 s 51072 99600 51128 99900 6 la_data_in[20]
port 130 nsew signal input
rlabel metal3 s 100 16128 400 16184 6 la_data_in[21]
port 131 nsew signal input
rlabel metal2 s 61824 99600 61880 99900 6 la_data_in[22]
port 132 nsew signal input
rlabel metal3 s 100 90384 400 90440 6 la_data_in[23]
port 133 nsew signal input
rlabel metal2 s 43344 99600 43400 99900 6 la_data_in[24]
port 134 nsew signal input
rlabel metal3 s 99600 24192 99900 24248 6 la_data_in[25]
port 135 nsew signal input
rlabel metal2 s 32592 100 32648 400 6 la_data_in[26]
port 136 nsew signal input
rlabel metal3 s 100 7392 400 7448 6 la_data_in[27]
port 137 nsew signal input
rlabel metal3 s 100 36624 400 36680 6 la_data_in[28]
port 138 nsew signal input
rlabel metal3 s 100 75936 400 75992 6 la_data_in[29]
port 139 nsew signal input
rlabel metal3 s 100 67536 400 67592 6 la_data_in[2]
port 140 nsew signal input
rlabel metal2 s 7728 99600 7784 99900 6 la_data_in[30]
port 141 nsew signal input
rlabel metal3 s 100 88704 400 88760 6 la_data_in[31]
port 142 nsew signal input
rlabel metal2 s 50400 99600 50456 99900 6 la_data_in[32]
port 143 nsew signal input
rlabel metal3 s 99600 85008 99900 85064 6 la_data_in[33]
port 144 nsew signal input
rlabel metal2 s 30912 99600 30968 99900 6 la_data_in[34]
port 145 nsew signal input
rlabel metal2 s 41664 99600 41720 99900 6 la_data_in[35]
port 146 nsew signal input
rlabel metal3 s 99600 54096 99900 54152 6 la_data_in[36]
port 147 nsew signal input
rlabel metal2 s 34608 100 34664 400 6 la_data_in[37]
port 148 nsew signal input
rlabel metal2 s 48048 100 48104 400 6 la_data_in[38]
port 149 nsew signal input
rlabel metal3 s 100 33600 400 33656 6 la_data_in[39]
port 150 nsew signal input
rlabel metal3 s 99600 61824 99900 61880 6 la_data_in[3]
port 151 nsew signal input
rlabel metal3 s 99600 1008 99900 1064 6 la_data_in[40]
port 152 nsew signal input
rlabel metal3 s 100 94416 400 94472 6 la_data_in[41]
port 153 nsew signal input
rlabel metal3 s 99600 72576 99900 72632 6 la_data_in[42]
port 154 nsew signal input
rlabel metal2 s 61488 100 61544 400 6 la_data_in[43]
port 155 nsew signal input
rlabel metal2 s 47376 99600 47432 99900 6 la_data_in[44]
port 156 nsew signal input
rlabel metal2 s 13440 99600 13496 99900 6 la_data_in[45]
port 157 nsew signal input
rlabel metal2 s 8736 99600 8792 99900 6 la_data_in[46]
port 158 nsew signal input
rlabel metal2 s 39648 99600 39704 99900 6 la_data_in[47]
port 159 nsew signal input
rlabel metal2 s 46032 100 46088 400 6 la_data_in[48]
port 160 nsew signal input
rlabel metal3 s 100 52080 400 52136 6 la_data_in[49]
port 161 nsew signal input
rlabel metal2 s 81984 99600 82040 99900 6 la_data_in[4]
port 162 nsew signal input
rlabel metal3 s 100 30576 400 30632 6 la_data_in[50]
port 163 nsew signal input
rlabel metal3 s 100 26880 400 26936 6 la_data_in[51]
port 164 nsew signal input
rlabel metal3 s 100 29904 400 29960 6 la_data_in[52]
port 165 nsew signal input
rlabel metal3 s 99600 3024 99900 3080 6 la_data_in[53]
port 166 nsew signal input
rlabel metal2 s 36624 100 36680 400 6 la_data_in[54]
port 167 nsew signal input
rlabel metal3 s 99600 90720 99900 90776 6 la_data_in[55]
port 168 nsew signal input
rlabel metal2 s 17136 100 17192 400 6 la_data_in[56]
port 169 nsew signal input
rlabel metal2 s 26208 99600 26264 99900 6 la_data_in[57]
port 170 nsew signal input
rlabel metal2 s 37632 99600 37688 99900 6 la_data_in[58]
port 171 nsew signal input
rlabel metal2 s 58800 100 58856 400 6 la_data_in[59]
port 172 nsew signal input
rlabel metal3 s 100 672 400 728 6 la_data_in[5]
port 173 nsew signal input
rlabel metal2 s 20160 100 20216 400 6 la_data_in[60]
port 174 nsew signal input
rlabel metal3 s 99600 35616 99900 35672 6 la_data_in[61]
port 175 nsew signal input
rlabel metal2 s 29904 99600 29960 99900 6 la_data_in[62]
port 176 nsew signal input
rlabel metal2 s 90720 99600 90776 99900 6 la_data_in[63]
port 177 nsew signal input
rlabel metal2 s 87024 99600 87080 99900 6 la_data_in[6]
port 178 nsew signal input
rlabel metal3 s 99600 53088 99900 53144 6 la_data_in[7]
port 179 nsew signal input
rlabel metal2 s 71232 100 71288 400 6 la_data_in[8]
port 180 nsew signal input
rlabel metal3 s 100 72240 400 72296 6 la_data_in[9]
port 181 nsew signal input
rlabel metal2 s 28224 99600 28280 99900 6 la_data_out[0]
port 182 nsew signal output
rlabel metal3 s 99600 41664 99900 41720 6 la_data_out[10]
port 183 nsew signal output
rlabel metal3 s 100 85680 400 85736 6 la_data_out[11]
port 184 nsew signal output
rlabel metal3 s 99600 55104 99900 55160 6 la_data_out[12]
port 185 nsew signal output
rlabel metal2 s 49392 99600 49448 99900 6 la_data_out[13]
port 186 nsew signal output
rlabel metal2 s 44352 99600 44408 99900 6 la_data_out[14]
port 187 nsew signal output
rlabel metal2 s 52752 100 52808 400 6 la_data_out[15]
port 188 nsew signal output
rlabel metal3 s 99600 46368 99900 46424 6 la_data_out[16]
port 189 nsew signal output
rlabel metal2 s 98448 99600 98504 99900 6 la_data_out[17]
port 190 nsew signal output
rlabel metal3 s 100 99120 400 99176 6 la_data_out[18]
port 191 nsew signal output
rlabel metal3 s 99600 62832 99900 62888 6 la_data_out[19]
port 192 nsew signal output
rlabel metal2 s 29904 100 29960 400 6 la_data_out[1]
port 193 nsew signal output
rlabel metal3 s 99600 28896 99900 28952 6 la_data_out[20]
port 194 nsew signal output
rlabel metal3 s 100 17136 400 17192 6 la_data_out[21]
port 195 nsew signal output
rlabel metal3 s 99600 12768 99900 12824 6 la_data_out[22]
port 196 nsew signal output
rlabel metal2 s 60816 99600 60872 99900 6 la_data_out[23]
port 197 nsew signal output
rlabel metal3 s 99600 79296 99900 79352 6 la_data_out[24]
port 198 nsew signal output
rlabel metal2 s 43344 100 43400 400 6 la_data_out[25]
port 199 nsew signal output
rlabel metal3 s 100 77952 400 78008 6 la_data_out[26]
port 200 nsew signal output
rlabel metal3 s 99600 45360 99900 45416 6 la_data_out[27]
port 201 nsew signal output
rlabel metal3 s 100 37632 400 37688 6 la_data_out[28]
port 202 nsew signal output
rlabel metal2 s 58800 99600 58856 99900 6 la_data_out[29]
port 203 nsew signal output
rlabel metal3 s 99600 18480 99900 18536 6 la_data_out[2]
port 204 nsew signal output
rlabel metal2 s 49056 100 49112 400 6 la_data_out[30]
port 205 nsew signal output
rlabel metal2 s 54096 99600 54152 99900 6 la_data_out[31]
port 206 nsew signal output
rlabel metal3 s 99600 80304 99900 80360 6 la_data_out[32]
port 207 nsew signal output
rlabel metal3 s 99600 38640 99900 38696 6 la_data_out[33]
port 208 nsew signal output
rlabel metal3 s 99600 2016 99900 2072 6 la_data_out[34]
port 209 nsew signal output
rlabel metal3 s 99600 13440 99900 13496 6 la_data_out[35]
port 210 nsew signal output
rlabel metal3 s 100 5712 400 5768 6 la_data_out[36]
port 211 nsew signal output
rlabel metal3 s 100 89712 400 89768 6 la_data_out[37]
port 212 nsew signal output
rlabel metal3 s 100 45024 400 45080 6 la_data_out[38]
port 213 nsew signal output
rlabel metal3 s 99600 84000 99900 84056 6 la_data_out[39]
port 214 nsew signal output
rlabel metal2 s 5712 100 5768 400 6 la_data_out[3]
port 215 nsew signal output
rlabel metal2 s 41328 100 41384 400 6 la_data_out[40]
port 216 nsew signal output
rlabel metal2 s 15456 99600 15512 99900 6 la_data_out[41]
port 217 nsew signal output
rlabel metal2 s 91392 100 91448 400 6 la_data_out[42]
port 218 nsew signal output
rlabel metal3 s 100 71232 400 71288 6 la_data_out[43]
port 219 nsew signal output
rlabel metal2 s 22848 100 22904 400 6 la_data_out[44]
port 220 nsew signal output
rlabel metal2 s 90384 100 90440 400 6 la_data_out[45]
port 221 nsew signal output
rlabel metal2 s 57120 99600 57176 99900 6 la_data_out[46]
port 222 nsew signal output
rlabel metal2 s 34944 99600 35000 99900 6 la_data_out[47]
port 223 nsew signal output
rlabel metal3 s 100 96432 400 96488 6 la_data_out[48]
port 224 nsew signal output
rlabel metal2 s 72576 99600 72632 99900 6 la_data_out[49]
port 225 nsew signal output
rlabel metal3 s 100 1680 400 1736 6 la_data_out[4]
port 226 nsew signal output
rlabel metal2 s 78288 99600 78344 99900 6 la_data_out[50]
port 227 nsew signal output
rlabel metal2 s 42672 99600 42728 99900 6 la_data_out[51]
port 228 nsew signal output
rlabel metal3 s 100 14448 400 14504 6 la_data_out[52]
port 229 nsew signal output
rlabel metal3 s 99600 58800 99900 58856 6 la_data_out[53]
port 230 nsew signal output
rlabel metal3 s 99600 68544 99900 68600 6 la_data_out[54]
port 231 nsew signal output
rlabel metal3 s 99600 88704 99900 88760 6 la_data_out[55]
port 232 nsew signal output
rlabel metal3 s 100 91392 400 91448 6 la_data_out[56]
port 233 nsew signal output
rlabel metal2 s 80976 99600 81032 99900 6 la_data_out[57]
port 234 nsew signal output
rlabel metal2 s 26880 100 26936 400 6 la_data_out[58]
port 235 nsew signal output
rlabel metal2 s 86688 100 86744 400 6 la_data_out[59]
port 236 nsew signal output
rlabel metal3 s 99600 6720 99900 6776 6 la_data_out[5]
port 237 nsew signal output
rlabel metal3 s 100 15120 400 15176 6 la_data_out[60]
port 238 nsew signal output
rlabel metal2 s 35616 99600 35672 99900 6 la_data_out[61]
port 239 nsew signal output
rlabel metal2 s 62496 100 62552 400 6 la_data_out[62]
port 240 nsew signal output
rlabel metal3 s 99600 47376 99900 47432 6 la_data_out[63]
port 241 nsew signal output
rlabel metal3 s 99600 37632 99900 37688 6 la_data_out[6]
port 242 nsew signal output
rlabel metal3 s 99600 70560 99900 70616 6 la_data_out[7]
port 243 nsew signal output
rlabel metal3 s 99600 56112 99900 56168 6 la_data_out[8]
port 244 nsew signal output
rlabel metal2 s 38640 99600 38696 99900 6 la_data_out[9]
port 245 nsew signal output
rlabel metal3 s 100 79968 400 80024 6 la_oenb[0]
port 246 nsew signal input
rlabel metal2 s 73248 100 73304 400 6 la_oenb[10]
port 247 nsew signal input
rlabel metal2 s 87696 100 87752 400 6 la_oenb[11]
port 248 nsew signal input
rlabel metal2 s 14448 100 14504 400 6 la_oenb[12]
port 249 nsew signal input
rlabel metal3 s 100 12432 400 12488 6 la_oenb[13]
port 250 nsew signal input
rlabel metal2 s 6720 99600 6776 99900 6 la_oenb[14]
port 251 nsew signal input
rlabel metal3 s 99600 8736 99900 8792 6 la_oenb[15]
port 252 nsew signal input
rlabel metal2 s 19488 99600 19544 99900 6 la_oenb[16]
port 253 nsew signal input
rlabel metal3 s 100 87696 400 87752 6 la_oenb[17]
port 254 nsew signal input
rlabel metal2 s 88032 99600 88088 99900 6 la_oenb[18]
port 255 nsew signal input
rlabel metal2 s 74256 99600 74312 99900 6 la_oenb[19]
port 256 nsew signal input
rlabel metal2 s 27888 100 27944 400 6 la_oenb[1]
port 257 nsew signal input
rlabel metal3 s 100 55776 400 55832 6 la_oenb[20]
port 258 nsew signal input
rlabel metal2 s 88704 100 88760 400 6 la_oenb[21]
port 259 nsew signal input
rlabel metal3 s 100 53760 400 53816 6 la_oenb[22]
port 260 nsew signal input
rlabel metal2 s 18144 100 18200 400 6 la_oenb[23]
port 261 nsew signal input
rlabel metal3 s 100 61488 400 61544 6 la_oenb[24]
port 262 nsew signal input
rlabel metal3 s 99600 94752 99900 94808 6 la_oenb[25]
port 263 nsew signal input
rlabel metal2 s 99456 99600 99512 99900 6 la_oenb[26]
port 264 nsew signal input
rlabel metal3 s 99600 86016 99900 86072 6 la_oenb[27]
port 265 nsew signal input
rlabel metal3 s 99600 81984 99900 82040 6 la_oenb[28]
port 266 nsew signal input
rlabel metal3 s 99600 80976 99900 81032 6 la_oenb[29]
port 267 nsew signal input
rlabel metal2 s 51072 100 51128 400 6 la_oenb[2]
port 268 nsew signal input
rlabel metal2 s 17472 99600 17528 99900 6 la_oenb[30]
port 269 nsew signal input
rlabel metal2 s 2688 100 2744 400 6 la_oenb[31]
port 270 nsew signal input
rlabel metal2 s 672 100 728 400 6 la_oenb[32]
port 271 nsew signal input
rlabel metal2 s 1008 99600 1064 99900 6 la_oenb[33]
port 272 nsew signal input
rlabel metal2 s 52080 100 52136 400 6 la_oenb[34]
port 273 nsew signal input
rlabel metal3 s 100 43344 400 43400 6 la_oenb[35]
port 274 nsew signal input
rlabel metal3 s 100 54768 400 54824 6 la_oenb[36]
port 275 nsew signal input
rlabel metal3 s 100 28896 400 28952 6 la_oenb[37]
port 276 nsew signal input
rlabel metal2 s 36624 99600 36680 99900 6 la_oenb[38]
port 277 nsew signal input
rlabel metal3 s 100 63504 400 63560 6 la_oenb[39]
port 278 nsew signal input
rlabel metal2 s 19152 100 19208 400 6 la_oenb[3]
port 279 nsew signal input
rlabel metal2 s 44352 100 44408 400 6 la_oenb[40]
port 280 nsew signal input
rlabel metal3 s 100 50064 400 50120 6 la_oenb[41]
port 281 nsew signal input
rlabel metal2 s 79968 100 80024 400 6 la_oenb[42]
port 282 nsew signal input
rlabel metal2 s 37632 100 37688 400 6 la_oenb[43]
port 283 nsew signal input
rlabel metal3 s 100 73248 400 73304 6 la_oenb[44]
port 284 nsew signal input
rlabel metal3 s 99600 48384 99900 48440 6 la_oenb[45]
port 285 nsew signal input
rlabel metal3 s 99600 66528 99900 66584 6 la_oenb[46]
port 286 nsew signal input
rlabel metal2 s 76944 100 77000 400 6 la_oenb[47]
port 287 nsew signal input
rlabel metal2 s 32928 99600 32984 99900 6 la_oenb[48]
port 288 nsew signal input
rlabel metal2 s 99120 100 99176 400 6 la_oenb[49]
port 289 nsew signal input
rlabel metal3 s 99600 63840 99900 63896 6 la_oenb[4]
port 290 nsew signal input
rlabel metal2 s 67536 99600 67592 99900 6 la_oenb[50]
port 291 nsew signal input
rlabel metal3 s 99600 51072 99900 51128 6 la_oenb[51]
port 292 nsew signal input
rlabel metal2 s 75936 100 75992 400 6 la_oenb[52]
port 293 nsew signal input
rlabel metal2 s 88704 99600 88760 99900 6 la_oenb[53]
port 294 nsew signal input
rlabel metal3 s 99600 9744 99900 9800 6 la_oenb[54]
port 295 nsew signal input
rlabel metal2 s 59808 99600 59864 99900 6 la_oenb[55]
port 296 nsew signal input
rlabel metal2 s 92400 100 92456 400 6 la_oenb[56]
port 297 nsew signal input
rlabel metal3 s 100 49056 400 49112 6 la_oenb[57]
port 298 nsew signal input
rlabel metal2 s 12432 100 12488 400 6 la_oenb[58]
port 299 nsew signal input
rlabel metal3 s 99600 50400 99900 50456 6 la_oenb[59]
port 300 nsew signal input
rlabel metal3 s 100 95424 400 95480 6 la_oenb[5]
port 301 nsew signal input
rlabel metal3 s 99600 65856 99900 65912 6 la_oenb[60]
port 302 nsew signal input
rlabel metal2 s 24864 100 24920 400 6 la_oenb[61]
port 303 nsew signal input
rlabel metal2 s 95424 100 95480 400 6 la_oenb[62]
port 304 nsew signal input
rlabel metal3 s 100 18144 400 18200 6 la_oenb[63]
port 305 nsew signal input
rlabel metal2 s 86016 99600 86072 99900 6 la_oenb[6]
port 306 nsew signal input
rlabel metal3 s 99600 76272 99900 76328 6 la_oenb[7]
port 307 nsew signal input
rlabel metal2 s 25200 99600 25256 99900 6 la_oenb[8]
port 308 nsew signal input
rlabel metal3 s 100 64512 400 64568 6 la_oenb[9]
port 309 nsew signal input
rlabel metal4 s 2224 1538 2384 98422 6 vdd
port 310 nsew power bidirectional
rlabel metal4 s 17584 1538 17744 98422 6 vdd
port 310 nsew power bidirectional
rlabel metal4 s 32944 1538 33104 98422 6 vdd
port 310 nsew power bidirectional
rlabel metal4 s 48304 1538 48464 98422 6 vdd
port 310 nsew power bidirectional
rlabel metal4 s 63664 1538 63824 98422 6 vdd
port 310 nsew power bidirectional
rlabel metal4 s 79024 1538 79184 98422 6 vdd
port 310 nsew power bidirectional
rlabel metal4 s 94384 1538 94544 98422 6 vdd
port 310 nsew power bidirectional
rlabel metal4 s 9904 1538 10064 98422 6 vss
port 311 nsew ground bidirectional
rlabel metal4 s 25264 1538 25424 98422 6 vss
port 311 nsew ground bidirectional
rlabel metal4 s 40624 1538 40784 98422 6 vss
port 311 nsew ground bidirectional
rlabel metal4 s 55984 1538 56144 98422 6 vss
port 311 nsew ground bidirectional
rlabel metal4 s 71344 1538 71504 98422 6 vss
port 311 nsew ground bidirectional
rlabel metal4 s 86704 1538 86864 98422 6 vss
port 311 nsew ground bidirectional
rlabel metal3 s 99600 17472 99900 17528 6 wb_clk_i
port 312 nsew signal input
rlabel metal2 s 18480 99600 18536 99900 6 wb_rst_i
port 313 nsew signal input
rlabel metal3 s 99600 34944 99900 35000 6 wbs_ack_o
port 314 nsew signal output
rlabel metal2 s 66528 99600 66584 99900 6 wbs_adr_i[0]
port 315 nsew signal input
rlabel metal2 s 45360 99600 45416 99900 6 wbs_adr_i[10]
port 316 nsew signal input
rlabel metal2 s 5712 99600 5768 99900 6 wbs_adr_i[11]
port 317 nsew signal input
rlabel metal2 s 8400 100 8456 400 6 wbs_adr_i[12]
port 318 nsew signal input
rlabel metal2 s 55776 100 55832 400 6 wbs_adr_i[13]
port 319 nsew signal input
rlabel metal3 s 99600 73584 99900 73640 6 wbs_adr_i[14]
port 320 nsew signal input
rlabel metal3 s 99600 67536 99900 67592 6 wbs_adr_i[15]
port 321 nsew signal input
rlabel metal2 s 63504 100 63560 400 6 wbs_adr_i[16]
port 322 nsew signal input
rlabel metal3 s 99600 59808 99900 59864 6 wbs_adr_i[17]
port 323 nsew signal input
rlabel metal3 s 99600 30912 99900 30968 6 wbs_adr_i[18]
port 324 nsew signal input
rlabel metal2 s 96432 100 96488 400 6 wbs_adr_i[19]
port 325 nsew signal input
rlabel metal3 s 100 6720 400 6776 6 wbs_adr_i[1]
port 326 nsew signal input
rlabel metal3 s 100 58800 400 58856 6 wbs_adr_i[20]
port 327 nsew signal input
rlabel metal2 s 56784 100 56840 400 6 wbs_adr_i[21]
port 328 nsew signal input
rlabel metal2 s 80976 100 81032 400 6 wbs_adr_i[22]
port 329 nsew signal input
rlabel metal3 s 99600 23184 99900 23240 6 wbs_adr_i[23]
port 330 nsew signal input
rlabel metal2 s 11760 99600 11816 99900 6 wbs_adr_i[24]
port 331 nsew signal input
rlabel metal2 s 54768 100 54824 400 6 wbs_adr_i[25]
port 332 nsew signal input
rlabel metal2 s 10416 100 10472 400 6 wbs_adr_i[26]
port 333 nsew signal input
rlabel metal2 s 33936 99600 33992 99900 6 wbs_adr_i[27]
port 334 nsew signal input
rlabel metal3 s 99600 58128 99900 58184 6 wbs_adr_i[28]
port 335 nsew signal input
rlabel metal3 s 99600 95760 99900 95816 6 wbs_adr_i[29]
port 336 nsew signal input
rlabel metal3 s 100 11424 400 11480 6 wbs_adr_i[2]
port 337 nsew signal input
rlabel metal3 s 100 39312 400 39368 6 wbs_adr_i[30]
port 338 nsew signal input
rlabel metal3 s 99600 42672 99900 42728 6 wbs_adr_i[31]
port 339 nsew signal input
rlabel metal2 s 77952 100 78008 400 6 wbs_adr_i[3]
port 340 nsew signal input
rlabel metal2 s 77280 99600 77336 99900 6 wbs_adr_i[4]
port 341 nsew signal input
rlabel metal2 s 75264 100 75320 400 6 wbs_adr_i[5]
port 342 nsew signal input
rlabel metal3 s 100 48048 400 48104 6 wbs_adr_i[6]
port 343 nsew signal input
rlabel metal2 s 4704 100 4760 400 6 wbs_adr_i[7]
port 344 nsew signal input
rlabel metal3 s 99600 0 99900 56 6 wbs_adr_i[8]
port 345 nsew signal input
rlabel metal3 s 99600 27216 99900 27272 6 wbs_adr_i[9]
port 346 nsew signal input
rlabel metal2 s 31920 99600 31976 99900 6 wbs_cyc_i
port 347 nsew signal input
rlabel metal3 s 99600 87024 99900 87080 6 wbs_dat_i[0]
port 348 nsew signal input
rlabel metal3 s 100 76944 400 77000 6 wbs_dat_i[10]
port 349 nsew signal input
rlabel metal3 s 100 84672 400 84728 6 wbs_dat_i[11]
port 350 nsew signal input
rlabel metal3 s 100 80976 400 81032 6 wbs_dat_i[12]
port 351 nsew signal input
rlabel metal2 s 3696 100 3752 400 6 wbs_dat_i[13]
port 352 nsew signal input
rlabel metal3 s 100 21168 400 21224 6 wbs_dat_i[14]
port 353 nsew signal input
rlabel metal3 s 99600 52080 99900 52136 6 wbs_dat_i[15]
port 354 nsew signal input
rlabel metal2 s 57792 100 57848 400 6 wbs_dat_i[16]
port 355 nsew signal input
rlabel metal2 s 68544 99600 68600 99900 6 wbs_dat_i[17]
port 356 nsew signal input
rlabel metal2 s 92736 99600 92792 99900 6 wbs_dat_i[18]
port 357 nsew signal input
rlabel metal2 s 5040 99600 5096 99900 6 wbs_dat_i[19]
port 358 nsew signal input
rlabel metal2 s 15120 100 15176 400 6 wbs_dat_i[1]
port 359 nsew signal input
rlabel metal3 s 100 24864 400 24920 6 wbs_dat_i[20]
port 360 nsew signal input
rlabel metal2 s 95760 99600 95816 99900 6 wbs_dat_i[21]
port 361 nsew signal input
rlabel metal3 s 100 59808 400 59864 6 wbs_dat_i[22]
port 362 nsew signal input
rlabel metal3 s 99600 78288 99900 78344 6 wbs_dat_i[23]
port 363 nsew signal input
rlabel metal3 s 99600 32928 99900 32984 6 wbs_dat_i[24]
port 364 nsew signal input
rlabel metal2 s 69216 100 69272 400 6 wbs_dat_i[25]
port 365 nsew signal input
rlabel metal2 s 82992 99600 83048 99900 6 wbs_dat_i[26]
port 366 nsew signal input
rlabel metal2 s 24192 99600 24248 99900 6 wbs_dat_i[27]
port 367 nsew signal input
rlabel metal2 s 31584 100 31640 400 6 wbs_dat_i[28]
port 368 nsew signal input
rlabel metal3 s 99600 60816 99900 60872 6 wbs_dat_i[29]
port 369 nsew signal input
rlabel metal2 s 81984 100 82040 400 6 wbs_dat_i[2]
port 370 nsew signal input
rlabel metal3 s 99600 29904 99900 29960 6 wbs_dat_i[30]
port 371 nsew signal input
rlabel metal3 s 100 52752 400 52808 6 wbs_dat_i[31]
port 372 nsew signal input
rlabel metal3 s 99600 4032 99900 4088 6 wbs_dat_i[3]
port 373 nsew signal input
rlabel metal2 s 16128 100 16184 400 6 wbs_dat_i[4]
port 374 nsew signal input
rlabel metal2 s 50064 100 50120 400 6 wbs_dat_i[5]
port 375 nsew signal input
rlabel metal3 s 99600 43344 99900 43400 6 wbs_dat_i[6]
port 376 nsew signal input
rlabel metal2 s 79296 99600 79352 99900 6 wbs_dat_i[7]
port 377 nsew signal input
rlabel metal3 s 99600 89712 99900 89768 6 wbs_dat_i[8]
port 378 nsew signal input
rlabel metal3 s 99600 5040 99900 5096 6 wbs_dat_i[9]
port 379 nsew signal input
rlabel metal3 s 100 20160 400 20216 6 wbs_dat_o[0]
port 380 nsew signal output
rlabel metal3 s 99600 57120 99900 57176 6 wbs_dat_o[10]
port 381 nsew signal output
rlabel metal2 s 1680 100 1736 400 6 wbs_dat_o[11]
port 382 nsew signal output
rlabel metal3 s 99600 91728 99900 91784 6 wbs_dat_o[12]
port 383 nsew signal output
rlabel metal2 s 75264 99600 75320 99900 6 wbs_dat_o[13]
port 384 nsew signal output
rlabel metal3 s 99600 11760 99900 11816 6 wbs_dat_o[14]
port 385 nsew signal output
rlabel metal2 s 71568 99600 71624 99900 6 wbs_dat_o[15]
port 386 nsew signal output
rlabel metal3 s 100 27888 400 27944 6 wbs_dat_o[16]
port 387 nsew signal output
rlabel metal3 s 100 31584 400 31640 6 wbs_dat_o[17]
port 388 nsew signal output
rlabel metal2 s 67536 100 67592 400 6 wbs_dat_o[18]
port 389 nsew signal output
rlabel metal2 s 0 100 56 400 6 wbs_dat_o[19]
port 390 nsew signal output
rlabel metal2 s 78960 100 79016 400 6 wbs_dat_o[1]
port 391 nsew signal output
rlabel metal3 s 100 47040 400 47096 6 wbs_dat_o[20]
port 392 nsew signal output
rlabel metal3 s 100 86688 400 86744 6 wbs_dat_o[21]
port 393 nsew signal output
rlabel metal2 s 27216 99600 27272 99900 6 wbs_dat_o[22]
port 394 nsew signal output
rlabel metal3 s 100 32592 400 32648 6 wbs_dat_o[23]
port 395 nsew signal output
rlabel metal2 s 21168 100 21224 400 6 wbs_dat_o[24]
port 396 nsew signal output
rlabel metal2 s 7392 100 7448 400 6 wbs_dat_o[25]
port 397 nsew signal output
rlabel metal2 s 52080 99600 52136 99900 6 wbs_dat_o[26]
port 398 nsew signal output
rlabel metal2 s 28896 99600 28952 99900 6 wbs_dat_o[27]
port 399 nsew signal output
rlabel metal2 s 53760 100 53816 400 6 wbs_dat_o[28]
port 400 nsew signal output
rlabel metal2 s 69552 99600 69608 99900 6 wbs_dat_o[29]
port 401 nsew signal output
rlabel metal3 s 99600 28224 99900 28280 6 wbs_dat_o[2]
port 402 nsew signal output
rlabel metal3 s 100 65520 400 65576 6 wbs_dat_o[30]
port 403 nsew signal output
rlabel metal3 s 99600 77280 99900 77336 6 wbs_dat_o[31]
port 404 nsew signal output
rlabel metal2 s 22176 100 22232 400 6 wbs_dat_o[3]
port 405 nsew signal output
rlabel metal2 s 38304 100 38360 400 6 wbs_dat_o[4]
port 406 nsew signal output
rlabel metal3 s 100 8400 400 8456 6 wbs_dat_o[5]
port 407 nsew signal output
rlabel metal3 s 99600 74256 99900 74312 6 wbs_dat_o[6]
port 408 nsew signal output
rlabel metal2 s 60480 100 60536 400 6 wbs_dat_o[7]
port 409 nsew signal output
rlabel metal2 s 65856 99600 65912 99900 6 wbs_dat_o[8]
port 410 nsew signal output
rlabel metal2 s 64848 99600 64904 99900 6 wbs_dat_o[9]
port 411 nsew signal output
rlabel metal3 s 100 92400 400 92456 6 wbs_sel_i[0]
port 412 nsew signal input
rlabel metal2 s 10752 99600 10808 99900 6 wbs_sel_i[1]
port 413 nsew signal input
rlabel metal2 s 72240 100 72296 400 6 wbs_sel_i[2]
port 414 nsew signal input
rlabel metal3 s 100 22176 400 22232 6 wbs_sel_i[3]
port 415 nsew signal input
rlabel metal3 s 100 82992 400 83048 6 wbs_stb_i
port 416 nsew signal input
rlabel metal3 s 99600 49392 99900 49448 6 wbs_we_i
port 417 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 100000 100000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 13785888
string GDS_FILE /home/videogamo/Work/gfmpw-0/caravel_hack_soc/openlane/caravel_hack_soc/runs/22_12_05_22_32/results/signoff/caravel_hack_soc.magic.gds
string GDS_START 455710
<< end >>

