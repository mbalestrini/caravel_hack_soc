* NGSPICE file created from caravel_hack_soc.ext - technology: gf180mcuC

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_1 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_2 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_2 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_1 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_2 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai31_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_1 A1 A2 A3 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_16 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux2_2 I0 I1 S Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_4 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_1 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_8 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_1 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_1 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_64 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_64 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_2 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__tiel abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__tiel ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_32 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_32 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or3_1 A1 A2 A3 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or2_1 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__filltie abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__filltie VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffq_1 D CLK Q VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffnq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffnq_1 D CLKN Q VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_1 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_1 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux4_1 I0 I1 I2 I3 S0 S1 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_1 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor2_1 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai22_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_1 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_4 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and2_1 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffq_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffq_2 D CLK Q VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_1 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_2 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_1 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__endcap abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__endcap VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__antenna abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__antenna I VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and3_1 A1 A2 A3 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai221_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai221_1 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_3 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_3 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_2 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_1 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xnor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xnor2_1 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_1 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor2_2 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_2 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_4 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_1 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai31_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_2 A1 A2 A3 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_2 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffnq_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffnq_2 D CLKN Q VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_2 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_1 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_2 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_2 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_1 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_4 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_2 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or4_1 A1 A2 A3 A4 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_2 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_4 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_2 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_4 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and4_2 A1 A2 A3 A4 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_4 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and2_2 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor3_2 A1 A2 A3 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and4_4 A1 A2 A3 A4 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_2 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_4 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai31_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_4 A1 A2 A3 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_4 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xnor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xnor3_1 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_4 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_4 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and4_1 A1 A2 A3 A4 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai32_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai32_2 A1 A2 A3 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_4 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_3 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_3 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor3_1 A1 A2 A3 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai221_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai221_4 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai221_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai221_2 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dlyb_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dlyb_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or2_2 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_4 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dlyd_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dlyd_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dlyc_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dlyc_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or4_2 A1 A2 A3 A4 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai222_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai222_2 A1 A2 B1 B2 C1 C2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai33_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai33_1 A1 A2 A3 B1 B2 B3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_3 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_3 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_4 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi222_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi222_1 A1 A2 B1 B2 C1 C2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__tieh abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__tieh Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai22_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_2 A1 A2 B1 B2 ZN VDD VSS
.ends

.subckt caravel_hack_soc io_in[0] io_in[10] io_in[11] io_in[12] io_in[13] io_in[14]
+ io_in[15] io_in[16] io_in[17] io_in[18] io_in[19] io_in[1] io_in[20] io_in[21] io_in[22]
+ io_in[23] io_in[24] io_in[25] io_in[26] io_in[27] io_in[28] io_in[29] io_in[2] io_in[30]
+ io_in[31] io_in[32] io_in[33] io_in[34] io_in[35] io_in[36] io_in[37] io_in[3] io_in[4]
+ io_in[5] io_in[6] io_in[7] io_in[8] io_in[9] io_oeb[0] io_oeb[10] io_oeb[11] io_oeb[12]
+ io_oeb[13] io_oeb[14] io_oeb[15] io_oeb[16] io_oeb[17] io_oeb[18] io_oeb[19] io_oeb[1]
+ io_oeb[20] io_oeb[21] io_oeb[22] io_oeb[23] io_oeb[24] io_oeb[25] io_oeb[26] io_oeb[27]
+ io_oeb[28] io_oeb[29] io_oeb[2] io_oeb[30] io_oeb[31] io_oeb[32] io_oeb[33] io_oeb[34]
+ io_oeb[35] io_oeb[36] io_oeb[37] io_oeb[3] io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7]
+ io_oeb[8] io_oeb[9] io_out[0] io_out[10] io_out[11] io_out[12] io_out[13] io_out[14]
+ io_out[15] io_out[16] io_out[17] io_out[18] io_out[19] io_out[1] io_out[20] io_out[21]
+ io_out[22] io_out[23] io_out[24] io_out[25] io_out[26] io_out[27] io_out[28] io_out[29]
+ io_out[2] io_out[30] io_out[31] io_out[32] io_out[33] io_out[34] io_out[35] io_out[36]
+ io_out[37] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7] io_out[8] io_out[9]
+ irq[0] irq[1] irq[2] la_data_in[0] la_data_in[10] la_data_in[11] la_data_in[12]
+ la_data_in[13] la_data_in[14] la_data_in[15] la_data_in[16] la_data_in[17] la_data_in[18]
+ la_data_in[19] la_data_in[1] la_data_in[20] la_data_in[21] la_data_in[22] la_data_in[23]
+ la_data_in[24] la_data_in[25] la_data_in[26] la_data_in[27] la_data_in[28] la_data_in[29]
+ la_data_in[2] la_data_in[30] la_data_in[31] la_data_in[32] la_data_in[33] la_data_in[34]
+ la_data_in[35] la_data_in[36] la_data_in[37] la_data_in[38] la_data_in[39] la_data_in[3]
+ la_data_in[40] la_data_in[41] la_data_in[42] la_data_in[43] la_data_in[44] la_data_in[45]
+ la_data_in[46] la_data_in[47] la_data_in[48] la_data_in[49] la_data_in[4] la_data_in[50]
+ la_data_in[51] la_data_in[52] la_data_in[53] la_data_in[54] la_data_in[55] la_data_in[56]
+ la_data_in[57] la_data_in[58] la_data_in[59] la_data_in[5] la_data_in[60] la_data_in[61]
+ la_data_in[62] la_data_in[63] la_data_in[6] la_data_in[7] la_data_in[8] la_data_in[9]
+ la_data_out[0] la_data_out[10] la_data_out[11] la_data_out[12] la_data_out[13] la_data_out[14]
+ la_data_out[15] la_data_out[16] la_data_out[17] la_data_out[18] la_data_out[19]
+ la_data_out[1] la_data_out[20] la_data_out[21] la_data_out[22] la_data_out[23] la_data_out[24]
+ la_data_out[25] la_data_out[26] la_data_out[27] la_data_out[28] la_data_out[29]
+ la_data_out[2] la_data_out[30] la_data_out[31] la_data_out[32] la_data_out[33] la_data_out[34]
+ la_data_out[35] la_data_out[36] la_data_out[37] la_data_out[38] la_data_out[39]
+ la_data_out[3] la_data_out[40] la_data_out[41] la_data_out[42] la_data_out[43] la_data_out[44]
+ la_data_out[45] la_data_out[46] la_data_out[47] la_data_out[48] la_data_out[49]
+ la_data_out[4] la_data_out[50] la_data_out[51] la_data_out[52] la_data_out[53] la_data_out[54]
+ la_data_out[55] la_data_out[56] la_data_out[57] la_data_out[58] la_data_out[59]
+ la_data_out[5] la_data_out[60] la_data_out[61] la_data_out[62] la_data_out[63] la_data_out[6]
+ la_data_out[7] la_data_out[8] la_data_out[9] la_oenb[0] la_oenb[10] la_oenb[11]
+ la_oenb[12] la_oenb[13] la_oenb[14] la_oenb[15] la_oenb[16] la_oenb[17] la_oenb[18]
+ la_oenb[19] la_oenb[1] la_oenb[20] la_oenb[21] la_oenb[22] la_oenb[23] la_oenb[24]
+ la_oenb[25] la_oenb[26] la_oenb[27] la_oenb[28] la_oenb[29] la_oenb[2] la_oenb[30]
+ la_oenb[31] la_oenb[32] la_oenb[33] la_oenb[34] la_oenb[35] la_oenb[36] la_oenb[37]
+ la_oenb[38] la_oenb[39] la_oenb[3] la_oenb[40] la_oenb[41] la_oenb[42] la_oenb[43]
+ la_oenb[44] la_oenb[45] la_oenb[46] la_oenb[47] la_oenb[48] la_oenb[49] la_oenb[4]
+ la_oenb[50] la_oenb[51] la_oenb[52] la_oenb[53] la_oenb[54] la_oenb[55] la_oenb[56]
+ la_oenb[57] la_oenb[58] la_oenb[59] la_oenb[5] la_oenb[60] la_oenb[61] la_oenb[62]
+ la_oenb[63] la_oenb[6] la_oenb[7] la_oenb[8] la_oenb[9] vdd vss wb_clk_i wb_rst_i
+ wbs_ack_o wbs_adr_i[0] wbs_adr_i[10] wbs_adr_i[11] wbs_adr_i[12] wbs_adr_i[13] wbs_adr_i[14]
+ wbs_adr_i[15] wbs_adr_i[16] wbs_adr_i[17] wbs_adr_i[18] wbs_adr_i[19] wbs_adr_i[1]
+ wbs_adr_i[20] wbs_adr_i[21] wbs_adr_i[22] wbs_adr_i[23] wbs_adr_i[24] wbs_adr_i[25]
+ wbs_adr_i[26] wbs_adr_i[27] wbs_adr_i[28] wbs_adr_i[29] wbs_adr_i[2] wbs_adr_i[30]
+ wbs_adr_i[31] wbs_adr_i[3] wbs_adr_i[4] wbs_adr_i[5] wbs_adr_i[6] wbs_adr_i[7] wbs_adr_i[8]
+ wbs_adr_i[9] wbs_cyc_i wbs_dat_i[0] wbs_dat_i[10] wbs_dat_i[11] wbs_dat_i[12] wbs_dat_i[13]
+ wbs_dat_i[14] wbs_dat_i[15] wbs_dat_i[16] wbs_dat_i[17] wbs_dat_i[18] wbs_dat_i[19]
+ wbs_dat_i[1] wbs_dat_i[20] wbs_dat_i[21] wbs_dat_i[22] wbs_dat_i[23] wbs_dat_i[24]
+ wbs_dat_i[25] wbs_dat_i[26] wbs_dat_i[27] wbs_dat_i[28] wbs_dat_i[29] wbs_dat_i[2]
+ wbs_dat_i[30] wbs_dat_i[31] wbs_dat_i[3] wbs_dat_i[4] wbs_dat_i[5] wbs_dat_i[6]
+ wbs_dat_i[7] wbs_dat_i[8] wbs_dat_i[9] wbs_dat_o[0] wbs_dat_o[10] wbs_dat_o[11]
+ wbs_dat_o[12] wbs_dat_o[13] wbs_dat_o[14] wbs_dat_o[15] wbs_dat_o[16] wbs_dat_o[17]
+ wbs_dat_o[18] wbs_dat_o[19] wbs_dat_o[1] wbs_dat_o[20] wbs_dat_o[21] wbs_dat_o[22]
+ wbs_dat_o[23] wbs_dat_o[24] wbs_dat_o[25] wbs_dat_o[26] wbs_dat_o[27] wbs_dat_o[28]
+ wbs_dat_o[29] wbs_dat_o[2] wbs_dat_o[30] wbs_dat_o[31] wbs_dat_o[3] wbs_dat_o[4]
+ wbs_dat_o[5] wbs_dat_o[6] wbs_dat_o[7] wbs_dat_o[8] wbs_dat_o[9] wbs_sel_i[0] wbs_sel_i[1]
+ wbs_sel_i[2] wbs_sel_i[3] wbs_stb_i wbs_we_i
XFILLER_41_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05903_ _01724_ _01728_ _01787_ _01789_ _01799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
X_09671_ _04639_ soc.rom_loader.current_address\[3\] _04647_ _04648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06883_ _02482_ _02492_ _02548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_05834_ _01732_ _01733_ _01729_ _01669_ _01734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_27_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08622_ _02149_ soc.spi_video_ram_1.write_fifo.fifo_mem\[30\]\[14\] _04011_ _04016_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_82_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_199_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05765_ _01662_ _01663_ _01661_ _01586_ _01668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_08553_ _03979_ _00466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_93_1615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_58_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07504_ _02903_ _03151_ _03152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_165_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08484_ _03942_ _00434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05696_ soc.cpu.AReg.data\[3\] soc.cpu.AReg.data\[2\] soc.cpu.AReg.data\[1\] _01603_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_1_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_161_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07435_ _03021_ soc.spi_video_ram_1.write_fifo.fifo_mem\[20\]\[27\] _03083_ _03084_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_52_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07366_ soc.spi_video_ram_1.output_buffer\[13\] _02676_ _03016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_52_1356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06317_ soc.spi_video_ram_1.fifo_in_address\[10\] _02173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_09105_ _02165_ soc.spi_video_ram_1.write_fifo.fifo_mem\[20\]\[22\] _04258_ _04283_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_109_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07297_ _02937_ _02946_ _02947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xcaravel_hack_soc_207 wbs_dat_o[15] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_178_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xcaravel_hack_soc_218 wbs_dat_o[26] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_09036_ soc.spi_video_ram_1.write_fifo.fifo_mem\[21\]\[28\] _02353_ _04221_ _04242_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06248_ _02126_ soc.spi_video_ram_1.write_fifo.fifo_mem\[18\]\[3\] _02120_ _02127_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_50_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_191_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_104_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06179_ soc.video_generator_1.h_count\[4\] _01836_ soc.video_generator_1.h_count\[6\]
+ _02068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_132_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_117_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_215_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_191_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_172_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_1430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09938_ soc.ram_encoder_0.input_bits_left\[3\] _04839_ _04841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_172_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_1463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_246_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_115_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_189_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09869_ soc.rom_encoder_0.request_data_out\[12\] _04742_ _04788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_85_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11900_ _00959_ clknet_leaf_296_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[3\]\[26\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_3246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_218_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11831_ _00890_ clknet_leaf_122_wb_clk_i soc.rom_encoder_0.input_buffer\[5\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_61_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1800 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_165_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1811 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1822 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_183_1242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1833 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1844 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11762_ _00823_ clknet_leaf_70_wb_clk_i soc.spi_video_ram_1.state_sram_clk_counter\[5\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_242_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1855 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1866 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_201_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10713_ _03443_ _05324_ _05337_ _01269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_13_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1877 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1888 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1899 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11693_ _00754_ clknet_leaf_130_wb_clk_i soc.spi_video_ram_1.fifo_in_data\[11\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_74_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10644_ _05300_ _01237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_10575_ _05259_ _05257_ _05260_ _01208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_10_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12314_ _01342_ clknet_leaf_155_wb_clk_i soc.ram_encoder_0.data_out\[9\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_202_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12245_ _01273_ clknet_leaf_273_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[29\]\[27\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12176_ _01204_ clknet_leaf_85_wb_clk_i soc.boot_loading_offset\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_9_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_237_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_1388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11127_ _00193_ clknet_leaf_192_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[14\]\[7\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_116_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11058_ _00124_ clknet_leaf_229_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[0\]\[25\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_5160 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5171 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_114_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5182 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_60_wb_clk_i clknet_5_12_0_wb_clk_i clknet_leaf_60_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_5193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10009_ soc.ram_encoder_0.request_data_out\[7\] soc.ram_encoder_0.data_out\[7\] _04889_
+ _04890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_4470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_149_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_184_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3780 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3791 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05550_ _01459_ _00011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_60_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_232_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_177_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05481_ _01395_ _01396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_18_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_92_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07220_ _02596_ _02871_ _02872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_34_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_73_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_242_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_220_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07151_ soc.spi_video_ram_1.write_fifo.fifo_mem\[0\]\[5\] soc.spi_video_ram_1.write_fifo.fifo_mem\[1\]\[5\]
+ soc.spi_video_ram_1.write_fifo.fifo_mem\[2\]\[5\] soc.spi_video_ram_1.write_fifo.fifo_mem\[3\]\[5\]
+ _02700_ _02647_ _02806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_06102_ soc.display_clks_before_active\[0\] _01903_ _01904_ _01995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_220_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07082_ _02726_ soc.spi_video_ram_1.write_fifo.fifo_mem\[4\]\[3\] _02739_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_106_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06033_ soc.video_generator_1.h_count\[1\] _01926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_160_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_234_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07984_ _02685_ _03623_ _02720_ _03624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09723_ _04678_ _04687_ _04688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_80_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06935_ _02570_ _02596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_67_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_228_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09654_ soc.rom_encoder_0.data_out\[14\] soc.rom_encoder_0.request_data_out\[14\]
+ _04632_ _04636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06866_ _01702_ _02535_ _02536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_83_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_242_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08605_ _02132_ soc.spi_video_ram_1.write_fifo.fifo_mem\[30\]\[6\] _04000_ _04007_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_05817_ soc.cpu.ALU.zy _01717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_06797_ _02443_ _02473_ _02474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09585_ _04590_ _04585_ _04591_ _00887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_58_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05748_ _01553_ soc.cpu.instruction\[3\] soc.cpu.AReg.data\[3\] _01592_ _01653_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_08536_ _03970_ _00458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_93_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_230_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_224_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05679_ _01560_ _01584_ _01586_ _01587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_50_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08467_ _03932_ _03933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_106_1508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07418_ _03065_ _03066_ _02958_ _03067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_08398_ soc.spi_video_ram_1.write_fifo.fifo_mem\[26\]\[27\] _02351_ _03865_ _03895_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_71_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_183_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07349_ _02941_ soc.spi_video_ram_1.write_fifo.fifo_mem\[23\]\[28\] _02690_ _02999_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_87_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10360_ soc.cpu.ALU.x\[14\] _05102_ _05120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_164_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09019_ _04233_ _00678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_124_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10291_ soc.rom_loader.current_address\[3\] _05076_ _05078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_105_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12030_ _01089_ clknet_leaf_67_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[5\]\[18\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_120_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_232_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3010 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_234_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_46_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3021 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3032 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3043 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3054 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xcaravel_hack_soc_94 io_oeb[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_3065 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3076 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3087 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3098 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_226_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11814_ _00873_ clknet_leaf_48_wb_clk_i soc.spi_video_ram_1.write_fifo.write_pointer\[1\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XTAP_1630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_183_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_214_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_159_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11745_ _00806_ clknet_leaf_75_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[4\]\[18\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1696 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_5_29_0_wb_clk_i clknet_4_14_0_wb_clk_i clknet_5_29_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_187_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_187_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11676_ _00737_ clknet_leaf_64_wb_clk_i soc.video_generator_1.v_count\[4\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_35_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_202_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10627_ soc.spi_video_ram_1.write_fifo.fifo_mem\[19\]\[12\] _04047_ _05289_ _05292_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_239_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_155_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10558_ soc.boot_loading_offset\[1\] _05246_ soc.boot_loading_offset\[2\] _05249_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_128_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_192_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10489_ _05172_ _05204_ _05205_ _01176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_29_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_1753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12228_ _01256_ clknet_leaf_16_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[29\]\[10\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_64_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12159_ _01187_ clknet_leaf_145_wb_clk_i soc.ram_encoder_0.address\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_64_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_111_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_204_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06720_ soc.spi_video_ram_1.write_fifo.fifo_mem\[14\]\[12\] _02242_ _02412_ _02416_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_65_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_224_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06651_ _02373_ _00171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_77_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_240_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05602_ _01507_ _01508_ _01509_ _01510_ _01469_ _01501_ _01511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_266_wb_clk_i clknet_5_7_0_wb_clk_i clknet_leaf_266_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_06582_ _02333_ _00142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09370_ soc.spi_video_ram_1.state_sram_clk_counter\[4\] _04439_ _04441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_212_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_206_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08321_ _03853_ _00360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05533_ _01405_ _01401_ _01442_ _01443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_32_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08252_ _02558_ _03809_ _03810_ _00334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_162_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05464_ _01379_ _01380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_138_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_203_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07203_ soc.spi_video_ram_1.write_fifo.fifo_mem\[4\]\[7\] soc.spi_video_ram_1.write_fifo.fifo_mem\[5\]\[7\]
+ soc.spi_video_ram_1.write_fifo.fifo_mem\[6\]\[7\] soc.spi_video_ram_1.write_fifo.fifo_mem\[7\]\[7\]
+ _02763_ _02838_ _02856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_165_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_159_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08183_ _03757_ _00318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_140_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_192_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07134_ _02678_ _02782_ _02789_ _02586_ _02790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_174_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07065_ soc.spi_video_ram_1.write_fifo.fifo_mem\[24\]\[2\] soc.spi_video_ram_1.write_fifo.fifo_mem\[25\]\[2\]
+ soc.spi_video_ram_1.write_fifo.fifo_mem\[26\]\[2\] soc.spi_video_ram_1.write_fifo.fifo_mem\[27\]\[2\]
+ _02689_ _02723_ _02724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_161_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06016_ _01883_ _01884_ _01909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_82_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_216_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_5907 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5918 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_47_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5929 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_102_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_210_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07967_ _02736_ _03607_ _03608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_116_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_151_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09706_ _04672_ soc.rom_encoder_0.request_address\[13\] _04617_ _04673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_28_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_216_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06918_ soc.spi_video_ram_1.write_fifo.fifo_mem\[12\]\[0\] soc.spi_video_ram_1.write_fifo.fifo_mem\[13\]\[0\]
+ soc.spi_video_ram_1.write_fifo.fifo_mem\[14\]\[0\] soc.spi_video_ram_1.write_fifo.fifo_mem\[15\]\[0\]
+ _02575_ _02578_ _02579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_229_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07898_ soc.spi_video_ram_1.write_fifo.fifo_mem\[15\]\[21\] _03541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_243_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09637_ soc.rom_encoder_0.data_out\[6\] soc.rom_encoder_0.request_data_out\[6\] _04621_
+ _04627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06849_ _02439_ soc.rom_encoder_0.output_bits_left\[2\] _02521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_245_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_227_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09568_ _04565_ _04574_ _04579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_231_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_208_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_149_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08519_ _03960_ _00451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_54_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_196_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09499_ _04534_ _00858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_51_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_157_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11530_ _00596_ clknet_leaf_278_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[23\]\[24\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_128_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11461_ _00527_ clknet_leaf_10_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[15\]\[13\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_128_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10412_ _02262_ soc.spi_video_ram_1.write_fifo.fifo_mem\[6\]\[22\] _05123_ _05148_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_11392_ _00458_ clknet_leaf_258_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[2\]\[2\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_178_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_193_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10343_ _01680_ _05103_ _05111_ _01125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_174_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10274_ soc.rom_loader.rom_request _04612_ soc.rom_loader.writing _05067_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_140_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_1355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_239_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12013_ _01072_ clknet_leaf_214_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[5\]\[1\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_79_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_171_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_235_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_246_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_206_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_222_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2150 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2161 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2172 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2183 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_221_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_14_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_206_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11728_ _00789_ clknet_leaf_227_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[4\]\[1\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_128_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_222_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_198_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11659_ _00720_ clknet_leaf_272_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[20\]\[27\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_156_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_200_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_174_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_196_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_1411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_233_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08870_ _04153_ _00609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_229_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07821_ _03047_ soc.spi_video_ram_1.write_fifo.fifo_mem\[14\]\[23\] _03465_ _02593_
+ _03466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_57_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_211_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07752_ _02893_ _03396_ _03397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_225_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06703_ _02404_ _00192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_65_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_1507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07683_ _02655_ _03305_ _03328_ _03329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_20_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09422_ soc.rom_encoder_0.request_data_out\[1\] _03767_ _04477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_25_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_241_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_198_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06634_ _02364_ _00163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_213_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_209_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09353_ soc.spi_video_ram_1.current_state\[3\] soc.spi_video_ram_1.current_state\[1\]
+ soc.spi_video_ram_1.current_state\[0\] soc.spi_video_ram_1.current_state\[2\] _04428_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
X_06565_ _02324_ _00134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_178_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08304_ _02145_ soc.spi_video_ram_1.write_fifo.fifo_mem\[1\]\[12\] _03842_ _03845_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_05516_ soc.spi_video_ram_1.initialized _01430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_06496_ _02285_ _00104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09284_ _04390_ _00786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_127_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08235_ soc.ram_encoder_0.output_buffer\[10\] _02563_ _03798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_105_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_193_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08166_ _02151_ soc.spi_video_ram_1.write_fifo.fifo_mem\[10\]\[15\] _03743_ _03749_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_134_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_238_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07117_ _02677_ _02606_ _02757_ _02773_ _02774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_08097_ soc.spi_video_ram_1.write_fifo.fifo_mem\[11\]\[26\] _02270_ _03679_ _03708_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_88_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07048_ _02706_ _02707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_122_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5704 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_62_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5715 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_134_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5726 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5737 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5748 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5759 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_134_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08999_ _04222_ _00669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_5_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_188_wb_clk_i clknet_5_29_0_wb_clk_i clknet_leaf_188_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_134_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_217_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_84_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_117_wb_clk_i clknet_5_26_0_wb_clk_i clknet_leaf_117_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_10961_ _00027_ clknet_leaf_10_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[18\]\[15\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_56_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_229_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_186_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_204_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_189_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10892_ _05434_ _01351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_203_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_245_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_197_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_200_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_223_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11513_ _00579_ clknet_leaf_195_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[23\]\[7\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_184_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_180_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12493_ net53 net52 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_8_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_201_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11444_ _00510_ clknet_leaf_231_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[30\]\[25\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_109_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_165_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_197_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11375_ _00441_ clknet_leaf_317_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[28\]\[14\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_10_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10326_ soc.rom_loader.wait_fall_clk soc.rom_loader.rom_request _00817_ _05101_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_113_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_180_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_152_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10257_ soc.spi_video_ram_1.fifo_in_address\[7\] _05045_ _05057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_3_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_230_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_1718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10188_ soc.hack_clock_0.counter\[0\] _05017_ _01064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_93_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_207_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_223_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_228_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_50_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_241_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06350_ _02180_ _02193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_128_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_187_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06281_ soc.spi_video_ram_1.fifo_in_data\[14\] _02149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_50_1432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_129_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08020_ _02736_ _03657_ _03658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_50_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_239_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_176_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_170_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09971_ _04863_ _04848_ _04864_ _01000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_170_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08922_ soc.spi_video_ram_1.write_fifo.fifo_mem\[22\]\[3\] _02397_ _04178_ _04182_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_48_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08853_ soc.spi_video_ram_1.write_fifo.fifo_mem\[25\]\[0\] _02310_ _04144_ _04145_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_131_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_242_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07804_ soc.spi_video_ram_1.write_fifo.fifo_mem\[0\]\[23\] soc.spi_video_ram_1.write_fifo.fifo_mem\[1\]\[23\]
+ soc.spi_video_ram_1.write_fifo.fifo_mem\[2\]\[23\] soc.spi_video_ram_1.write_fifo.fifo_mem\[3\]\[23\]
+ _02680_ _02838_ _03449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
Xclkbuf_leaf_281_wb_clk_i clknet_5_4_0_wb_clk_i clknet_leaf_281_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_61_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08784_ soc.spi_video_ram_1.write_fifo.fifo_mem\[24\]\[28\] _02353_ _04075_ _04106_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_05996_ _01880_ _01888_ _01855_ _01889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_66_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_210_wb_clk_i clknet_5_20_0_wb_clk_i clknet_leaf_210_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_38_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07735_ soc.spi_video_ram_1.write_fifo.fifo_mem\[18\]\[15\] soc.spi_video_ram_1.write_fifo.fifo_mem\[19\]\[15\]
+ _02597_ _03380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_2908 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2919 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_246_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07666_ soc.spi_video_ram_1.write_fifo.fifo_mem\[15\]\[14\] _03312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_168_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_164_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09405_ _02542_ _04461_ _04462_ _04463_ _00835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_164_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06617_ _02354_ _00156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_81_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_240_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07597_ _02618_ _03243_ _03244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_179_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09336_ _02262_ soc.spi_video_ram_1.write_fifo.fifo_mem\[4\]\[22\] _04394_ _04419_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_107_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06548_ _02116_ _02313_ _02314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_142_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_205_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_166_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09267_ _02256_ soc.spi_video_ram_1.write_fifo.fifo_mem\[9\]\[19\] _04359_ _04382_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_103_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06479_ soc.spi_video_ram_1.write_fifo.fifo_mem\[16\]\[28\] _02274_ _02216_ _02275_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_138_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08218_ soc.ram_encoder_0.output_buffer\[6\] _02563_ _03785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09198_ _00011_ _01652_ _04344_ _00746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_135_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08149_ _02134_ soc.spi_video_ram_1.write_fifo.fifo_mem\[10\]\[7\] _03732_ _03740_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_194_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_179_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11160_ _00226_ clknet_leaf_92_wb_clk_i soc.rom_encoder_0.output_buffer\[3\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_49_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_6202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10111_ soc.ram_encoder_0.request_data_out\[7\] _04930_ _04959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_161_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11091_ _00157_ clknet_leaf_177_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[12\]\[0\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_6235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10042_ soc.ram_encoder_0.request_address\[7\] soc.ram_encoder_0.address\[7\] _04900_
+ _04907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_231_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4800 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_195_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4811 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_5567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4822 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4833 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_236_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4844 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4855 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4866 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4877 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4888 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4899 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11993_ _01052_ clknet_leaf_117_wb_clk_i soc.ram_data_out\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_1_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_205_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_147_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10944_ soc.spi_video_ram_1.write_fifo.fifo_mem\[8\]\[28\] soc.spi_video_ram_1.fifo_in_address\[12\]
+ _05430_ _05461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_229_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_232_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10875_ _01779_ _05221_ _05411_ _05424_ _01344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_16_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_38_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xclkbuf_leaf_85_wb_clk_i clknet_5_14_0_wb_clk_i clknet_leaf_85_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XPHY_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_185_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_157_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_14_wb_clk_i clknet_5_2_0_wb_clk_i clknet_leaf_14_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_138_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_5 soc.rom_encoder_0.data_out\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11427_ _00493_ clknet_leaf_179_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[30\]\[8\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_158_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_236_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_152_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11358_ _00424_ clknet_leaf_293_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[27\]\[26\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_158_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_193_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10309_ soc.rom_loader.current_address\[9\] _05088_ _05090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_234_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11289_ _00355_ clknet_leaf_0_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[1\]\[15\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_140_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_1583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_171_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_239_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05850_ _01722_ _01738_ _01747_ _01749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_43_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_212_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05781_ _01558_ soc.cpu.ALU.x\[6\] _01683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_187_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07520_ _02597_ soc.spi_video_ram_1.write_fifo.fifo_mem\[12\]\[26\] _02943_ _03168_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_63_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_165_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_78_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07451_ _02767_ _03094_ _03099_ _02970_ _03100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_63_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_222_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_1319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06402_ soc.spi_video_ram_1.fifo_in_data\[3\] _02223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_50_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07382_ _03027_ _03028_ _03030_ _02691_ _02588_ _03031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_37_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09121_ _01394_ _01429_ _01438_ _04291_ _04292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_176_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_163_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_06333_ _02184_ _00042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_143_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_148_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06264_ _02137_ _00020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09052_ _04243_ _04252_ _04253_ _00691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_191_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_198_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08003_ _02768_ _03641_ _03642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_102_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06195_ _01476_ _02081_ _02082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_144_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_opt_5_0_wb_clk_i clknet_5_31_0_wb_clk_i clknet_opt_5_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_190_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_171_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_1_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_143_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09954_ soc.ram_encoder_0.input_buffer\[2\] _04853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_83_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08905_ _04171_ _00626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09885_ _02436_ _02454_ soc.rom_encoder_0.current_state\[2\] _04800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4107 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4118 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_218_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4129 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08836_ _04063_ _04124_ _04135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_100_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_211_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08767_ _04097_ _00562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2705 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05979_ soc.video_generator_1.v_count\[9\] soc.video_generator_1.v_count\[1\] _01850_
+ _01871_ _01872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_122_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2716 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2727 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07718_ soc.spi_video_ram_1.write_fifo.fifo_mem\[9\]\[24\] _03364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_2738 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2749 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08698_ _04058_ _00532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_214_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07649_ _02601_ _03294_ _03295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_241_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_198_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_246_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10660_ _05308_ _01245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_16_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_224_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09319_ _04410_ _00801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_167_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10591_ soc.gpio_i_stored\[1\] _05268_ _02053_ _05271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_22_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12330_ _01358_ clknet_leaf_200_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[8\]\[9\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_202_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_194_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_12261_ _01289_ clknet_leaf_315_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[31\]\[14\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_110_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_208_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_123_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11212_ _00278_ clknet_leaf_254_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[11\]\[22\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_134_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12192_ _01220_ clknet_leaf_143_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[19\]\[3\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_150_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6010 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput53 net53 io_oeb[19] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_11143_ _00209_ clknet_leaf_284_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[14\]\[23\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_6021 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput64 net64 io_out[16] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_96_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_6032 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput75 net75 io_out[28] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_235_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_89_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6043 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_132_wb_clk_i clknet_5_24_0_wb_clk_i clknet_leaf_132_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_6054 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6065 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11074_ _00140_ clknet_leaf_7_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[13\]\[12\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_6076 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_118_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6087 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_49_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6098 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10025_ soc.ram_encoder_0.request_data_out\[15\] soc.ram_encoder_0.data_out\[15\]
+ _04889_ _04898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_88_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_237_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_49_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_149_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3940 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4696 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3951 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3962 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3973 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11976_ _01035_ clknet_leaf_153_wb_clk_i soc.ram_encoder_0.request_address\[13\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3984 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3995 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10927_ _05452_ _01368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_204_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_242_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_220_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10858_ soc.ram_encoder_0.data_out\[3\] _05416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_34_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_158_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10789_ _02213_ soc.spi_video_ram_1.write_fifo.fifo_mem\[7\]\[0\] _05378_ _05379_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XPHY_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_200_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_184_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_199_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_201_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_86_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06951_ _02572_ _02612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_80_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_214_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05902_ _01791_ _01795_ _01797_ _01798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_09670_ _04639_ _04646_ _04647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_132_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06882_ _02547_ _00228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_223_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08621_ _04015_ _00498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_227_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05833_ _01725_ _01727_ _01733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_167_1408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08552_ _02140_ soc.spi_video_ram_1.write_fifo.fifo_mem\[2\]\[10\] _03978_ _03979_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_05764_ _01595_ _01666_ _01667_ soc.cpu.PC.in\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_70_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07503_ soc.spi_video_ram_1.write_fifo.fifo_mem\[23\]\[26\] _03151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_78_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_39_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08483_ _02134_ soc.spi_video_ram_1.write_fifo.fifo_mem\[28\]\[7\] _03934_ _03942_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_223_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05695_ net78 _01564_ _01576_ _01577_ _01602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_22_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07434_ _03054_ soc.spi_video_ram_1.write_fifo.fifo_mem\[21\]\[27\] _03083_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_168_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_23_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07365_ _02624_ _02882_ _03015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_206_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_241_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09104_ _04282_ _00714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_176_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06316_ _02172_ _00037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_164_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07296_ _02707_ _02938_ _02945_ _02910_ _02946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_11_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xcaravel_hack_soc_208 wbs_dat_o[16] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xcaravel_hack_soc_219 wbs_dat_o[27] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_09035_ _04241_ _00686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_164_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06247_ soc.spi_video_ram_1.fifo_in_data\[3\] _02126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_102_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_176_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06178_ soc.video_generator_1.h_count\[4\] _01836_ soc.video_generator_1.h_count\[6\]
+ _02067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_105_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09937_ _02480_ _04839_ _04840_ _00990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_172_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_232_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_217_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_131_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_154_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09868_ _01395_ _04787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_219_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_133_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08819_ _04126_ _00585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_86_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09799_ _02111_ _02456_ _04731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_3236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_189_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11830_ _00889_ clknet_leaf_123_wb_clk_i soc.rom_encoder_0.input_buffer\[4\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_2_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1801 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1823 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1834 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11761_ _00822_ clknet_leaf_70_wb_clk_i soc.spi_video_ram_1.state_sram_clk_counter\[4\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_57_1246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_144_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_41_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_199_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_187_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1856 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10712_ soc.spi_video_ram_1.fifo_in_address\[7\] _05325_ _05337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_1867 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_5_19_0_wb_clk_i clknet_4_9_0_wb_clk_i clknet_5_19_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XTAP_1878 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_202_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1889 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11692_ _00753_ clknet_leaf_132_wb_clk_i soc.spi_video_ram_1.fifo_in_data\[10\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_70_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10643_ soc.spi_video_ram_1.write_fifo.fifo_mem\[19\]\[20\] soc.spi_video_ram_1.fifo_in_address\[4\]
+ _05277_ _05300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_201_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10574_ _01452_ _05260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_166_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12313_ _01341_ clknet_leaf_155_wb_clk_i soc.ram_encoder_0.data_out\[8\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_182_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_68_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12244_ _01272_ clknet_leaf_294_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[29\]\[26\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_leaf_313_wb_clk_i clknet_5_1_0_wb_clk_i clknet_leaf_313_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_6_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_155_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12175_ _01203_ clknet_leaf_85_wb_clk_i soc.boot_loading_offset\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_29_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_96_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11126_ _00192_ clknet_leaf_202_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[14\]\[6\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_110_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_218_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5150 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11057_ _00123_ clknet_leaf_296_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[0\]\[24\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_114_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5161 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5172 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_231_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5183 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10008_ _04879_ _04889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_209_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_236_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_149_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_209_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3770 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3781 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3792 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11959_ _01018_ clknet_leaf_114_wb_clk_i soc.ram_encoder_0.request_data_out\[12\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_33_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_205_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_1414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_209_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_199_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05480_ _01378_ _01395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_189_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_20_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_207_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_186_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_201_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07150_ _02596_ _02804_ _02640_ _02805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_146_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_158_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_185_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06101_ soc.display_clks_before_active\[0\] _01994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_9_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07081_ soc.spi_video_ram_1.write_fifo.fifo_mem\[0\]\[3\] soc.spi_video_ram_1.write_fifo.fifo_mem\[1\]\[3\]
+ soc.spi_video_ram_1.write_fifo.fifo_mem\[2\]\[3\] soc.spi_video_ram_1.write_fifo.fifo_mem\[3\]\[3\]
+ _02713_ _02737_ _02738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_103_1480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06032_ _01901_ _01905_ _01925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_86_1442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_236_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07983_ soc.spi_video_ram_1.write_fifo.fifo_mem\[4\]\[18\] soc.spi_video_ram_1.write_fifo.fifo_mem\[5\]\[18\]
+ soc.spi_video_ram_1.write_fifo.fifo_mem\[6\]\[18\] soc.spi_video_ram_1.write_fifo.fifo_mem\[7\]\[18\]
+ _02717_ _02682_ _03623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_113_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09722_ _04681_ _04682_ _04686_ _04687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_80_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06934_ _02589_ _02594_ _02595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_151_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09653_ _04635_ _00911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06865_ _01670_ soc.cpu.ALU.x\[15\] _02535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_27_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_28_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08604_ _04006_ _00490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_110_1440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05816_ _01702_ _01715_ _01716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_167_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09584_ net7 _04586_ _04553_ _04591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_3_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06796_ soc.rom_encoder_0.output_buffer\[19\] _02463_ _02464_ soc.rom_encoder_0.request_data_out\[15\]
+ _02473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08535_ _02124_ soc.spi_video_ram_1.write_fifo.fifo_mem\[2\]\[2\] _03967_ _03970_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_05747_ _01615_ _01651_ _01652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_169_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_242_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08466_ _03931_ _02214_ _03932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05678_ _01585_ _01586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_195_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07417_ _02696_ soc.spi_video_ram_1.write_fifo.fifo_mem\[12\]\[27\] _03066_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_52_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08397_ _03894_ _00395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_104_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07348_ _02613_ soc.spi_video_ram_1.write_fifo.fifo_mem\[22\]\[28\] _02998_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_104_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_192_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07279_ _02569_ _02929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_164_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09018_ soc.spi_video_ram_1.write_fifo.fifo_mem\[21\]\[19\] _02341_ _04221_ _04233_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_136_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10290_ soc.rom_loader.current_address\[3\] _05076_ _05077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_117_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_215_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3000 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3011 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3022 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3033 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_218_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3044 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3055 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xcaravel_hack_soc_95 io_oeb[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_73_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3066 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3077 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_234_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11813_ _00872_ clknet_leaf_60_wb_clk_i soc.spi_video_ram_1.write_fifo.write_pointer\[0\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3088 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3099 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_183_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11744_ _00805_ clknet_leaf_67_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[4\]\[17\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_226_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1697 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_230_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11675_ _00736_ clknet_leaf_129_wb_clk_i soc.video_generator_1.v_count\[3\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_169_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_168_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10626_ _05291_ _01228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_128_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10557_ _05248_ _01202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_6_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10488_ soc.cpu.PC.in\[10\] _05188_ _05201_ _05205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_155_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12227_ _01255_ clknet_leaf_255_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[29\]\[9\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_64_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_237_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_97_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_135_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12158_ _01186_ clknet_leaf_145_wb_clk_i soc.ram_encoder_0.address\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_150_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11109_ _00175_ clknet_leaf_28_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[12\]\[18\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_4_12_0_wb_clk_i clknet_3_6_0_wb_clk_i clknet_4_12_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_190_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12089_ soc.cpu.PC.in\[12\] net89 soc.cpu.AReg.data\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_238_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_168_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_237_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06650_ _02149_ soc.spi_video_ram_1.write_fifo.fifo_mem\[12\]\[14\] _02368_ _02373_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_77_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05601_ soc.spi_video_ram_1.output_buffer\[16\] _01510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_06581_ soc.spi_video_ram_1.write_fifo.fifo_mem\[13\]\[14\] _02246_ _02328_ _02333_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_220_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_224_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08320_ _02161_ soc.spi_video_ram_1.write_fifo.fifo_mem\[1\]\[20\] _03830_ _03853_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_162_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05532_ _01405_ _01401_ _01441_ _01398_ _01442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_244_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_177_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_205_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08251_ soc.ram_encoder_0.output_buffer\[14\] _02555_ _03810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_33_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05463_ _01378_ _01379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_4
XFILLER_127_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_193_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_242_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_220_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07202_ soc.spi_video_ram_1.write_fifo.fifo_mem\[8\]\[7\] soc.spi_video_ram_1.write_fifo.fifo_mem\[9\]\[7\]
+ soc.spi_video_ram_1.write_fifo.fifo_mem\[10\]\[7\] soc.spi_video_ram_1.write_fifo.fifo_mem\[11\]\[7\]
+ _02680_ _02722_ _02855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
Xclkbuf_leaf_235_wb_clk_i clknet_5_16_0_wb_clk_i clknet_leaf_235_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_197_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08182_ _02167_ soc.spi_video_ram_1.write_fifo.fifo_mem\[10\]\[23\] _03731_ _03757_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_146_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07133_ _02693_ _02786_ _02787_ _02788_ _02643_ _02789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_119_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07064_ _02722_ _02723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_118_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06015_ _01900_ _01906_ _01907_ _01908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_5908 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_134_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5919 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07966_ soc.spi_video_ram_1.write_fifo.fifo_mem\[24\]\[19\] soc.spi_video_ram_1.write_fifo.fifo_mem\[25\]\[19\]
+ soc.spi_video_ram_1.write_fifo.fifo_mem\[26\]\[19\] soc.spi_video_ram_1.write_fifo.fifo_mem\[27\]\[19\]
+ _02713_ _02737_ _03607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_09705_ soc.cpu.PC.REG.data\[13\] soc.rom_loader.current_address\[13\] _04638_ _04672_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06917_ _02577_ _02578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_68_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_228_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07897_ _03535_ _03536_ _03539_ _02691_ _02929_ _03540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_83_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09636_ _04626_ _00903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_28_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06848_ _02519_ _02520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_167_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_216_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09567_ _04576_ _04578_ _00882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06779_ _02456_ _02457_ _02458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_71_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_230_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_243_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_145_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08518_ _02169_ soc.spi_video_ram_1.write_fifo.fifo_mem\[28\]\[24\] _03933_ _03960_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_12_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09498_ _02252_ soc.cpu.AReg.data\[1\] _04339_ _04534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_180_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_227_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08449_ _03922_ _00419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_212_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_196_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_184_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_183_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11460_ _00526_ clknet_leaf_308_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[15\]\[12\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_137_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_177_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_149_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10411_ _05147_ _01157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_11391_ _00457_ clknet_leaf_212_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[2\]\[1\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_197_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_158_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10342_ soc.cpu.ALU.x\[5\] _05109_ _05111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_87_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_109_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_30_1282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_3_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_69_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10273_ _03714_ _05066_ _01100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_3_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12012_ _01071_ clknet_leaf_212_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[5\]\[0\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_152_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_61_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xclkbuf_leaf_39_wb_clk_i clknet_5_3_0_wb_clk_i clknet_leaf_39_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_82_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_1468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_43_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_232_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_246_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_219_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_210_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_185_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_235_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2140 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2151 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_1722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_206_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2162 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2173 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2184 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11727_ _00788_ clknet_leaf_214_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[4\]\[0\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_124_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_202_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_243_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11658_ _00719_ clknet_leaf_287_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[20\]\[26\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_30_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_190_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_11_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10609_ _05282_ _01220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_11589_ _00655_ clknet_leaf_242_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[22\]\[25\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_122_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_9_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_135_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07820_ _02613_ _03464_ _03465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_111_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_245_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07751_ soc.spi_video_ram_1.write_fifo.fifo_mem\[29\]\[15\] _03396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_22_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_5_1_0_wb_clk_i clknet_4_0_0_wb_clk_i clknet_5_1_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_65_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06702_ soc.spi_video_ram_1.write_fifo.fifo_mem\[14\]\[6\] _02403_ _02391_ _02404_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_77_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07682_ _02655_ _03318_ _03327_ _03328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_37_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_231_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09421_ _04473_ _04475_ _04476_ _00838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06633_ _02132_ soc.spi_video_ram_1.write_fifo.fifo_mem\[12\]\[6\] _02357_ _02364_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_92_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_212_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_225_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09352_ _04427_ _00817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_80_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06564_ soc.spi_video_ram_1.write_fifo.fifo_mem\[13\]\[6\] _02229_ _02317_ _02324_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_08303_ _03844_ _00351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_100_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05515_ _01428_ _01417_ _01429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09283_ _02272_ soc.spi_video_ram_1.write_fifo.fifo_mem\[9\]\[27\] _04359_ _04390_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_142_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06495_ _02130_ soc.spi_video_ram_1.write_fifo.fifo_mem\[0\]\[5\] _02279_ _02285_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_08234_ soc.ram_encoder_0.output_buffer\[6\] _03781_ _03789_ soc.ram_encoder_0.request_data_out\[2\]
+ _03796_ _03797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_20_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_140_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08165_ _03748_ _00309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_88_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_222_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_134_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_147_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07116_ _02760_ _02762_ _02766_ _02772_ _02568_ _02773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_175_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08096_ _03707_ _00281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_161_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07047_ _00002_ _02706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_6406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_216_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_138_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5705 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5716 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_114_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_5727 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5738 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5749 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_197_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08998_ soc.spi_video_ram_1.write_fifo.fifo_mem\[21\]\[10\] _02411_ _04221_ _04222_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_75_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_235_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07949_ _02768_ _03590_ _03591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_151_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_229_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_229_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_21_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10960_ _00026_ clknet_leaf_4_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[18\]\[14\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_90_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_217_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09619_ _01379_ _04611_ _04615_ _04616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_182_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10891_ soc.spi_video_ram_1.write_fifo.fifo_mem\[8\]\[2\] soc.spi_video_ram_1.fifo_in_data\[2\]
+ _05431_ _05434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_231_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xclkbuf_leaf_157_wb_clk_i clknet_5_27_0_wb_clk_i clknet_leaf_157_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_38_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_70_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_19_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_238_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_12_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11512_ _00578_ clknet_leaf_247_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[23\]\[6\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12492_ net53 net51 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_240_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_200_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11443_ _00509_ clknet_leaf_300_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[30\]\[24\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_123_1483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11374_ _00440_ clknet_leaf_311_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[28\]\[13\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_124_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_193_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10325_ net45 _05100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_98_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_238_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10256_ _03504_ _05044_ _05056_ _01093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_45_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_78_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10187_ _01380_ _05016_ _05017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_113_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_227_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_207_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_206_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_06280_ _02148_ _00025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_198_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_200_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_190_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_235_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09970_ soc.ram_encoder_0.input_buffer\[3\] _04849_ _04248_ _04864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_171_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_217_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08921_ _04181_ _00632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_139_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08852_ _04143_ _04144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_07803_ _03430_ _03438_ _03447_ _02567_ _03448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_112_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_217_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08783_ _04105_ _00570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05995_ _01881_ _01878_ _01887_ _01868_ _01888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XFILLER_72_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07734_ _03379_ _00247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_66_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2909 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_241_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07665_ _03306_ _03307_ _03310_ _02690_ _02569_ _03311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_198_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_183_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_213_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09404_ soc.rom_encoder_0.request_address\[4\] _02543_ _04463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_25_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06616_ soc.spi_video_ram_1.write_fifo.fifo_mem\[13\]\[28\] _02353_ _02316_ _02354_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xclkbuf_leaf_250_wb_clk_i clknet_5_17_0_wb_clk_i clknet_leaf_250_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_80_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07596_ _02984_ _03239_ _03242_ _03243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_197_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09335_ _04418_ _00809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_94_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_200_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06547_ soc.spi_video_ram_1.write_fifo.write_pointer\[4\] _02312_ _02313_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_244_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09266_ _04381_ _00777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06478_ soc.spi_video_ram_1.fifo_in_address\[12\] _02274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_08217_ soc.ram_encoder_0.request_address\[5\] _02506_ _03781_ soc.ram_encoder_0.output_buffer\[2\]
+ _03784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_193_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09197_ soc.spi_video_ram_1.fifo_in_data\[3\] _04341_ _04344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_217_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08148_ _03739_ _00301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_106_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_194_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08079_ soc.spi_video_ram_1.write_fifo.fifo_mem\[11\]\[17\] _02337_ _03691_ _03699_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_122_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10110_ _04952_ _04958_ _01044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_6214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_175_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_6225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11090_ _00156_ clknet_leaf_282_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[13\]\[28\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_6236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10041_ _04906_ _01028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_6269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_130_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_209_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4801 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_212_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4812 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4823 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4834 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_188_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4845 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4856 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4867 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4878 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11992_ _01051_ clknet_leaf_118_wb_clk_i soc.ram_data_out\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_75_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4889 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_112_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_186_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10943_ _05460_ _01376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_72_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10874_ soc.ram_encoder_0.data_out\[11\] _05424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_147_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_73_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_242_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_223_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_129_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_184_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_199_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_61_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_201_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_177_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11426_ _00492_ clknet_leaf_193_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[30\]\[7\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_6 net15 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_54_wb_clk_i clknet_5_24_0_wb_clk_i clknet_leaf_54_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_158_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11357_ _00423_ clknet_leaf_231_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[27\]\[25\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_141_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10308_ soc.rom_loader.current_address\[9\] _05088_ _05089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_113_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11288_ _00354_ clknet_leaf_317_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[1\]\[14\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_3_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10239_ soc.spi_video_ram_1.fifo_in_data\[14\] _05045_ _05048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_79_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05780_ _01586_ _01682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_35_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_223_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_228_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07450_ _03095_ _03096_ _03098_ _02958_ _02642_ _03099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_62_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_211_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06401_ _02222_ _00072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_241_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07381_ _02926_ soc.spi_video_ram_1.write_fifo.fifo_mem\[20\]\[11\] _03029_ _03030_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_52_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09120_ _04290_ _02673_ _01434_ _01419_ _04291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_06332_ _02122_ soc.spi_video_ram_1.write_fifo.fifo_mem\[17\]\[1\] _02182_ _02184_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_176_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09051_ soc.spi_video_ram_1.write_fifo.read_pointer\[3\] _04251_ _04253_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_175_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06263_ _02136_ soc.spi_video_ram_1.write_fifo.fifo_mem\[18\]\[8\] _02120_ _02137_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_08002_ soc.spi_video_ram_1.write_fifo.fifo_mem\[0\]\[17\] soc.spi_video_ram_1.write_fifo.fifo_mem\[1\]\[17\]
+ soc.spi_video_ram_1.write_fifo.fifo_mem\[2\]\[17\] soc.spi_video_ram_1.write_fifo.fifo_mem\[3\]\[17\]
+ _02769_ _02758_ _03641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_191_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06194_ _01516_ _01522_ _01524_ _01471_ _02081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_239_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_219_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_176_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09953_ _04851_ _04848_ _04852_ _00994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_103_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_48_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08904_ soc.spi_video_ram_1.write_fifo.fifo_mem\[25\]\[25\] _04069_ _04143_ _04171_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_170_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09884_ _04787_ _04799_ _00978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4108 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_246_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_213_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4119 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08835_ _03554_ _04124_ _04134_ _00593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_3407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08766_ soc.spi_video_ram_1.write_fifo.fifo_mem\[24\]\[19\] _02341_ _04087_ _04097_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_3429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05978_ soc.boot_loading_offset\[1\] _01871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_57_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2706 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2717 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07717_ _02703_ soc.spi_video_ram_1.write_fifo.fifo_mem\[11\]\[24\] _02646_ _03363_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_2728 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_187_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08697_ soc.spi_video_ram_1.write_fifo.fifo_mem\[15\]\[18\] _02339_ _04043_ _04058_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_2739 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_199_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_198_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07648_ _03289_ _03290_ _03293_ _02581_ _03294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_246_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_26_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_81_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07579_ _03139_ _03225_ _03226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_15_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_201_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_146_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09318_ _02244_ soc.spi_video_ram_1.write_fifo.fifo_mem\[4\]\[13\] _04406_ _04410_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_51_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_220_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10590_ net15 _05270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_139_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09249_ _04372_ _00769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_127_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12260_ _01288_ clknet_leaf_314_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[31\]\[13\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_120_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_194_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11211_ _00277_ clknet_leaf_282_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[11\]\[21\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_103_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_12191_ _01219_ clknet_leaf_137_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[19\]\[2\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_123_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_218_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_6000 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11142_ _00208_ clknet_leaf_268_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[14\]\[22\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_6011 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput54 net54 io_oeb[22] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_6022 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput65 net65 io_out[17] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_6033 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput76 net76 io_out[29] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_6044 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6055 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11073_ _00139_ clknet_leaf_38_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[13\]\[11\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_231_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6066 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6077 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6088 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10024_ _04897_ _01020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_7_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6099 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_23_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_236_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_114_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3930 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3941 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3952 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4697 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_101_wb_clk_i clknet_5_14_0_wb_clk_i clknet_leaf_101_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_205_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3963 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11975_ _01034_ clknet_leaf_168_wb_clk_i soc.ram_encoder_0.request_address\[12\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3974 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_229_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3985 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3996 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_232_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10926_ soc.spi_video_ram_1.write_fifo.fifo_mem\[8\]\[19\] soc.spi_video_ram_1.fifo_in_address\[3\]
+ _05442_ _05452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_166_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10857_ _01632_ _05222_ _05412_ _05415_ _01335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_73_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10788_ _05377_ _05378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XPHY_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_185_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_160_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_121_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_242_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_157_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11409_ _00475_ clknet_leaf_74_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[2\]\[19\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_236_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_193_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06950_ _02583_ _02610_ _02586_ _02611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_98_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_171_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_239_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_228_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05901_ _01796_ _01797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_67_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06881_ soc.rom_encoder_0.output_buffer\[1\] _02542_ _02543_ soc.rom_encoder_0.request_address\[0\]
+ _02547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_08620_ _02147_ soc.spi_video_ram_1.write_fifo.fifo_mem\[30\]\[13\] _04011_ _04015_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_05832_ _01662_ _01691_ _01723_ _01732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_95_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08551_ _03965_ _03978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_05763_ _01553_ soc.cpu.instruction\[4\] soc.cpu.AReg.data\[4\] _01592_ _01667_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_82_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07502_ _02744_ soc.spi_video_ram_1.write_fifo.fifo_mem\[20\]\[26\] _03149_ _02927_
+ _03150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_78_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08482_ _03941_ _00433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05694_ net38 _01601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_63_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07433_ _03068_ _03074_ _03081_ _02655_ _03082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_56_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_210_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07364_ _01419_ _02917_ _03013_ _02677_ _03014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_148_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_221_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09103_ _02163_ soc.spi_video_ram_1.write_fifo.fifo_mem\[20\]\[21\] _04258_ _04282_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06315_ _02171_ soc.spi_video_ram_1.write_fifo.fifo_mem\[18\]\[25\] _02119_ _02172_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_104_1426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07295_ _02939_ _02940_ _02942_ _02944_ _02706_ _02945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_136_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09034_ soc.spi_video_ram_1.write_fifo.fifo_mem\[21\]\[27\] _02351_ _04221_ _04241_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xcaravel_hack_soc_209 wbs_dat_o[17] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_06246_ _02125_ _00014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_163_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06177_ soc.spi_video_ram_1.sram_sio_oe net57 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_190_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_219_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_191_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_132_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09936_ soc.ram_encoder_0.input_bits_left\[2\] _04838_ _04840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_63_1465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_232_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_218_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09867_ _04752_ _04786_ _00974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_1517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08818_ _02147_ soc.spi_video_ram_1.write_fifo.fifo_mem\[23\]\[13\] _04117_ _04126_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_3215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_234_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09798_ soc.rom_encoder_0.initializing_step\[1\] _02459_ _04729_ _04730_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_27_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08749_ _04088_ _00553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1802 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_214_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1813 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11760_ _00821_ clknet_leaf_70_wb_clk_i soc.spi_video_ram_1.state_sram_clk_counter\[3\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffnq_2
XTAP_1824 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_226_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1835 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_241_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1846 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_198_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10711_ _03494_ _05324_ _05336_ _01268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_1857 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_183_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1868 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11691_ _00752_ clknet_leaf_141_wb_clk_i soc.spi_video_ram_1.fifo_in_data\[9\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_144_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1879 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_224_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10642_ _05299_ _01236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_41_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_167_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_220_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_139_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10573_ soc.hack_wait_clocks\[1\] _05259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_6_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_70_1469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_194_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12312_ _01340_ clknet_leaf_155_wb_clk_i soc.ram_encoder_0.data_out\[7\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_33_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12243_ _01271_ clknet_leaf_290_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[29\]\[25\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_170_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_237_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_155_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_12174_ _01202_ clknet_leaf_126_wb_clk_i soc.boot_loading_offset\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_68_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_190_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_1357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11125_ _00191_ clknet_leaf_221_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[14\]\[5\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_123_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_5140 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11056_ _00122_ clknet_leaf_242_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[0\]\[23\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_5151 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_237_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5162 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5173 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10007_ _04888_ _01012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_49_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5184 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_49_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_133_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3760 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3771 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3782 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_233_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3793 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11958_ _01017_ clknet_leaf_118_wb_clk_i soc.ram_encoder_0.request_data_out\[11\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_45_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10909_ _05443_ _01359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_220_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11889_ _00948_ clknet_leaf_320_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[3\]\[15\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_60_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06100_ soc.video_generator_1.h_count\[3\] soc.video_generator_1.h_count\[2\] _01993_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_34_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_199_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07080_ _02636_ _02737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_66_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_218_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_201_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_173_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06031_ _01923_ _01924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_12_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_172_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_86_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_114_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_25_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07982_ _02768_ _03621_ _03622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_138_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_141_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09721_ _04683_ _02549_ _04684_ _04685_ _04686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_132_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06933_ soc.spi_video_ram_1.write_fifo.fifo_mem\[0\]\[0\] soc.spi_video_ram_1.write_fifo.fifo_mem\[1\]\[0\]
+ soc.spi_video_ram_1.write_fifo.fifo_mem\[2\]\[0\] soc.spi_video_ram_1.write_fifo.fifo_mem\[3\]\[0\]
+ _02591_ _02593_ _02594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_214_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09652_ soc.rom_encoder_0.data_out\[13\] soc.rom_encoder_0.request_data_out\[13\]
+ _04632_ _04635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06864_ _01705_ _02533_ _02534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_80_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_227_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_216_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08603_ _02130_ soc.spi_video_ram_1.write_fifo.fifo_mem\[30\]\[5\] _04000_ _04006_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_05815_ _01670_ soc.cpu.ALU.x\[8\] _01715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09583_ soc.rom_encoder_0.input_buffer\[2\] _04590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_06795_ _02453_ _02471_ _02472_ _01381_ _00216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_23_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08534_ _03969_ _00457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_70_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05746_ _01586_ _01648_ _01650_ _01651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_223_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08465_ _02115_ _02312_ _03862_ _03931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_169_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05677_ soc.cpu.ALU.f _01585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_23_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_243_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_196_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07416_ _02971_ soc.spi_video_ram_1.write_fifo.fifo_mem\[13\]\[27\] _03065_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_225_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_211_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08396_ soc.spi_video_ram_1.write_fifo.fifo_mem\[26\]\[26\] _02270_ _03865_ _03894_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_10_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07347_ _02691_ _02993_ _02996_ _02582_ _02997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_195_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07278_ _02926_ soc.spi_video_ram_1.write_fifo.fifo_mem\[9\]\[10\] _02927_ _02928_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_100_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_164_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09017_ _04232_ _00677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06229_ soc.ram_encoder_0.toggled_sram_sck _02112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_191_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_191_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_232_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09919_ soc.rom_encoder_0.initializing_step\[3\] _04825_ _04826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_8_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_219_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3001 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3012 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3023 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3034 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3045 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_189_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_46_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3056 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xcaravel_hack_soc_96 io_oeb[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_2322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3067 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3078 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3089 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11812_ _00871_ clknet_leaf_63_wb_clk_i soc.spi_video_ram_1.initialized vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_215_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_199_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11743_ _00804_ clknet_leaf_74_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[4\]\[16\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_18_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_202_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1698 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11674_ _00735_ clknet_leaf_128_wb_clk_i soc.video_generator_1.v_count\[2\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_70_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10625_ soc.spi_video_ram_1.write_fifo.fifo_mem\[19\]\[11\] _02414_ _05289_ _05291_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_204_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10556_ soc.boot_loading_offset\[1\] _05246_ _05247_ _05248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_155_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_196_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_182_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_185_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10487_ soc.cpu.PC.REG.data\[10\] _05203_ _05204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_6_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_170_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12226_ _01254_ clknet_leaf_177_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[29\]\[8\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_194_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_29_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_190_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12157_ _01185_ clknet_leaf_147_wb_clk_i soc.ram_encoder_0.address\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_29_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11108_ _00174_ clknet_leaf_21_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[12\]\[17\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_81_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12088_ soc.cpu.PC.in\[11\] net84 soc.cpu.AReg.data\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_231_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11039_ _00105_ clknet_leaf_247_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[0\]\[6\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_209_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05600_ soc.spi_video_ram_1.output_buffer\[18\] _01509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_18_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06580_ _02332_ _00141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_75_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_205_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05531_ soc.spi_video_ram_1.write_fifo.write_pointer\[1\] _01405_ _01441_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_162_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_221_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_178_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08250_ soc.ram_encoder_0.output_buffer\[10\] _03781_ _03789_ soc.ram_encoder_0.request_data_out\[6\]
+ _03808_ _03809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_05462_ net18 _01378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_222_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_207_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07201_ soc.spi_video_ram_1.write_fifo.fifo_mem\[12\]\[7\] soc.spi_video_ram_1.write_fifo.fifo_mem\[13\]\[7\]
+ soc.spi_video_ram_1.write_fifo.fifo_mem\[14\]\[7\] soc.spi_video_ram_1.write_fifo.fifo_mem\[15\]\[7\]
+ _02680_ _02838_ _02854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_177_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08181_ _03756_ _00317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_158_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_9_wb_clk_i clknet_5_3_0_wb_clk_i clknet_leaf_9_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_146_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07132_ _02726_ soc.spi_video_ram_1.write_fifo.fifo_mem\[14\]\[4\] _02770_ _02788_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_9_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07063_ _02646_ _02722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_179_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06014_ _01894_ _01899_ _01893_ _01907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_114_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5909 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_173_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07965_ _03599_ _03601_ _03603_ _03605_ _02710_ _03606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_114_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09704_ _04671_ _00926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_60_1446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06916_ _02576_ _02577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_60_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07896_ _02752_ soc.spi_video_ram_1.write_fifo.fifo_mem\[8\]\[21\] _03538_ _03539_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_95_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09635_ soc.rom_encoder_0.data_out\[5\] soc.rom_encoder_0.request_data_out\[5\] _04621_
+ _04626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06847_ _02454_ _02515_ _02463_ _02519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_244_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09566_ soc.rom_encoder_0.current_state\[2\] _04577_ _04578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06778_ _02435_ _02433_ _02457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_58_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_70_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05729_ _01617_ _01626_ _01634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_08517_ _03959_ _00450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_24_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09497_ _04533_ _00857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_180_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08448_ soc.spi_video_ram_1.write_fifo.fifo_mem\[27\]\[21\] _02260_ _03898_ _03922_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_141_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_208_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_71_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08379_ _03885_ _00386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_123_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10410_ _02260_ soc.spi_video_ram_1.write_fifo.fifo_mem\[6\]\[21\] _05123_ _05147_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_139_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_221_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11390_ _00456_ clknet_leaf_207_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[2\]\[0\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_109_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_87_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10341_ _01666_ _05103_ _05110_ _01124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_178_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_238_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_139_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10272_ soc.rom_loader.rom_request _05065_ _04611_ _05066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_65_1313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_1482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12011_ _01070_ clknet_leaf_113_wb_clk_i soc.hack_clock_0.counter\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_105_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_79_wb_clk_i clknet_5_10_0_wb_clk_i clknet_leaf_79_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_62_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_234_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2130 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_185_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2141 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2152 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2163 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2174 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2185 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_203_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_226_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11726_ _00787_ clknet_leaf_274_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[9\]\[28\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_230_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11657_ _00718_ clknet_leaf_235_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[20\]\[25\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_141_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10608_ soc.spi_video_ram_1.write_fifo.fifo_mem\[19\]\[3\] _02397_ _05278_ _05282_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_11588_ _00654_ clknet_leaf_277_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[22\]\[24\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_102_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_183_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10539_ _05239_ _01193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_7_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_155_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_237_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_12209_ _01237_ clknet_leaf_51_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[19\]\[20\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_97_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_238_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07750_ _02752_ soc.spi_video_ram_1.write_fifo.fifo_mem\[30\]\[15\] _03394_ _02827_
+ _03395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_133_1282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06701_ soc.spi_video_ram_1.fifo_in_data\[6\] _02403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_168_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07681_ _02706_ _03319_ _03326_ _02600_ _03327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_237_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_226_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09420_ soc.rom_encoder_0.output_buffer\[8\] _02542_ _04476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06632_ _02363_ _00162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_52_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09351_ _04426_ _01378_ _04427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06563_ _02323_ _00133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_244_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_205_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08302_ _02143_ soc.spi_video_ram_1.write_fifo.fifo_mem\[1\]\[11\] _03842_ _03844_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_05514_ soc.spi_video_ram_1.current_state\[3\] _01428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_09282_ _04389_ _00785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_90_1439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06494_ _02284_ _00103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08233_ soc.ram_encoder_0.request_address\[9\] _02505_ _03796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_220_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08164_ _02149_ soc.spi_video_ram_1.write_fifo.fifo_mem\[10\]\[14\] _03743_ _03748_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_181_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07115_ _02768_ _02771_ _02772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_146_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08095_ soc.spi_video_ram_1.write_fifo.fifo_mem\[11\]\[25\] _02268_ _03679_ _03707_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_162_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_118_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07046_ _02704_ soc.spi_video_ram_1.write_fifo.fifo_mem\[7\]\[2\] _02691_ _02705_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_115_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_88_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_6418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_192_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5706 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_47_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5717 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5728 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_130_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_216_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5739 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_134_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08997_ _04209_ _04221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_75_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07948_ soc.spi_video_ram_1.write_fifo.fifo_mem\[16\]\[20\] soc.spi_video_ram_1.write_fifo.fifo_mem\[17\]\[20\]
+ soc.spi_video_ram_1.write_fifo.fifo_mem\[18\]\[20\] soc.spi_video_ram_1.write_fifo.fifo_mem\[19\]\[20\]
+ _02764_ _02723_ _03590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_21_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_228_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_55_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07879_ _02677_ _02918_ _03499_ _03522_ _03523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_44_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_216_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09618_ _04614_ _04615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_147_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10890_ _05433_ _01350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_243_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09549_ _04243_ _04250_ _04251_ _00879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_24_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_240_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_227_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_212_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_145_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11511_ _00577_ clknet_leaf_213_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[23\]\[5\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_145_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_197_wb_clk_i clknet_5_25_0_wb_clk_i clknet_leaf_197_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_196_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12491_ net53 net50 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_180_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xclkbuf_leaf_126_wb_clk_i clknet_5_14_0_wb_clk_i clknet_leaf_126_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_11442_ _00508_ clknet_leaf_232_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[30\]\[23\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_171_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11373_ _00439_ clknet_leaf_6_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[28\]\[12\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_158_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10324_ _05071_ _05099_ _01117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_3_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_125_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_171_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10255_ soc.spi_video_ram_1.fifo_in_address\[6\] _05045_ _05056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_124_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_152_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_234_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10186_ soc.hack_clock_0.counter\[1\] _05012_ _05015_ _05016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_171_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_232_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_120_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_187_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_219_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_208_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_235_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_61_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_245_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_163_1242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_231_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_202_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11709_ _00770_ clknet_leaf_42_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[9\]\[11\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_124_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_89_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_226_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_196_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08920_ soc.spi_video_ram_1.write_fifo.fifo_mem\[22\]\[2\] _02395_ _04178_ _04181_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_130_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_174_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08851_ _04142_ _04143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_58_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_217_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07802_ _02901_ _03439_ _03446_ _02970_ _03447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_57_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05994_ _01883_ _01884_ _01877_ _01886_ _01887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
X_08782_ soc.spi_video_ram_1.write_fifo.fifo_mem\[24\]\[27\] _02351_ _04075_ _04105_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_22_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07733_ soc.spi_video_ram_1.output_buffer\[9\] _02882_ _03378_ _03379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_26_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_187_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_246_1317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_168_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07664_ _02590_ soc.spi_video_ram_1.write_fifo.fifo_mem\[8\]\[14\] _03309_ _03310_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_53_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_65_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09403_ soc.rom_encoder_0.output_buffer\[5\] _02541_ _04462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_225_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_164_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06615_ soc.spi_video_ram_1.fifo_in_address\[12\] _02353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_168_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07595_ _02689_ soc.spi_video_ram_1.write_fifo.fifo_mem\[20\]\[25\] _03241_ _02742_
+ _03242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_34_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_222_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_181_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09334_ _02260_ soc.spi_video_ram_1.write_fifo.fifo_mem\[4\]\[21\] _04394_ _04418_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06546_ _01403_ _02312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_142_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_194_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_221_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_290_wb_clk_i clknet_5_5_0_wb_clk_i clknet_leaf_290_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_06477_ _02273_ _00097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09265_ _02254_ soc.spi_video_ram_1.write_fifo.fifo_mem\[9\]\[18\] _04359_ _04381_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_178_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08216_ _02556_ _03782_ _03783_ _00325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_14_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09196_ _00011_ _01632_ _04343_ _00745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_222_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08147_ _02132_ soc.spi_video_ram_1.write_fifo.fifo_mem\[10\]\[6\] _03732_ _03739_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_147_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_200_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08078_ _03698_ _00272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_136_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_235_1722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07029_ _02644_ _02688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_1_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10040_ soc.ram_encoder_0.request_address\[6\] soc.ram_encoder_0.address\[6\] _04900_
+ _04906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_6259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4802 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4813 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4824 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_102_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_233_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4835 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_1171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_229_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4846 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4857 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4868 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4879 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11991_ _01050_ clknet_leaf_118_wb_clk_i soc.ram_data_out\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_17_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_60_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_217_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10942_ soc.spi_video_ram_1.write_fifo.fifo_mem\[8\]\[27\] soc.spi_video_ram_1.fifo_in_address\[11\]
+ _05430_ _05460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_44_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_231_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10873_ _01767_ _05221_ _05411_ _05423_ _01343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_38_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xclkbuf_leaf_307_wb_clk_i clknet_5_3_0_wb_clk_i clknet_leaf_307_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XPHY_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_101_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_213_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_125_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_240_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_200_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11425_ _00491_ clknet_leaf_210_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[30\]\[6\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_126_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_7 net23 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_193_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11356_ _00422_ clknet_leaf_298_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[27\]\[24\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10307_ _05071_ _05087_ _05088_ _01111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_4_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_112_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_193_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11287_ _00353_ clknet_leaf_319_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[1\]\[13\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10238_ _03225_ _05044_ _05047_ _01084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_80_1427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_leaf_23_wb_clk_i clknet_5_8_0_wb_clk_i clknet_leaf_23_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_10169_ _04919_ _05001_ _05002_ _03714_ _01060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_94_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_187_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_212_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_207_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06400_ soc.spi_video_ram_1.write_fifo.fifo_mem\[16\]\[2\] _02221_ _02217_ _02222_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_206_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_204_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07380_ _02919_ soc.spi_video_ram_1.write_fifo.fifo_mem\[21\]\[11\] _03029_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_96_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_194_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06331_ _02183_ _00041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_128_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_203_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_198_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09050_ soc.spi_video_ram_1.write_fifo.read_pointer\[3\] _04251_ _04252_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_176_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06262_ soc.spi_video_ram_1.fifo_in_data\[8\] _02136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_15_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_176_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08001_ _03577_ _03639_ _03579_ _03640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_190_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06193_ _02073_ _02079_ _02080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_129_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_219_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_237_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09952_ net2 _04849_ _04601_ _04852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_171_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08903_ _04170_ _00625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_106_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09883_ _01553_ _04741_ _04798_ _04799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4109 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08834_ _04061_ _04124_ _04134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_230_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08765_ _04096_ _00561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05977_ _01860_ _01866_ _01863_ _01870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_100_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2707 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07716_ _02903_ soc.spi_video_ram_1.write_fifo.fifo_mem\[10\]\[24\] _03362_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_2718 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2729 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08696_ _04057_ _00531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_57_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_183_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_213_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_14_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07647_ _02783_ soc.spi_video_ram_1.write_fifo.fifo_mem\[20\]\[14\] _03292_ _02741_
+ _03293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_96_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_246_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_228_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07578_ soc.spi_video_ram_1.write_fifo.fifo_mem\[5\]\[13\] _03225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_181_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09317_ _04409_ _00800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_181_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06529_ _02302_ _00120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_21_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09248_ _02237_ soc.spi_video_ram_1.write_fifo.fifo_mem\[9\]\[10\] _04365_ _04372_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_90_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_193_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_182_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_108_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09179_ _01849_ _01939_ _02034_ _04325_ _04332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_147_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11210_ _00276_ clknet_leaf_52_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[11\]\[20\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12190_ _01218_ clknet_leaf_219_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[19\]\[1\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_190_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11141_ _00207_ clknet_leaf_282_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[14\]\[21\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_6001 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_107_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6012 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_194_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xoutput55 net55 io_oeb[23] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_81_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6023 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput66 net66 io_out[18] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_62_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6034 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput77 net77 io_out[34] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_150_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11072_ _00138_ clknet_leaf_16_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[13\]\[10\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_6045 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6056 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_1_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_6067 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6078 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10023_ soc.ram_encoder_0.request_data_out\[14\] soc.ram_encoder_0.data_out\[14\]
+ _04889_ _04897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_76_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6089 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_4654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3920 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3931 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3942 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4698 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3953 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11974_ _01033_ clknet_leaf_153_wb_clk_i soc.ram_encoder_0.request_address\[11\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3964 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3975 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3986 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3997 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10925_ _05451_ _01367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_244_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_189_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_225_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_147_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_141_wb_clk_i clknet_5_25_0_wb_clk_i clknet_leaf_141_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_207_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10856_ soc.ram_encoder_0.data_out\[2\] _05415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_60_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_232_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_129_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_73_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10787_ _01445_ _04392_ _05377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XPHY_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_199_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_160_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_201_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_158_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_117_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11408_ _00474_ clknet_leaf_77_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[2\]\[18\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_114_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11339_ _00405_ clknet_leaf_186_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[27\]\[7\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_136_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05900_ _01782_ _01785_ _01796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_234_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06880_ _02546_ _00227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_6590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_95_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05831_ _01724_ _01728_ _01730_ _01731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_67_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_43_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05762_ _01654_ _01665_ _01666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_3_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08550_ _03977_ _00465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_242_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_229_wb_clk_i clknet_5_16_0_wb_clk_i clknet_leaf_229_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_78_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_236_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07501_ _02903_ _03148_ _03149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_63_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05693_ _01598_ _01599_ _01600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08481_ _02132_ soc.spi_video_ram_1.write_fifo.fifo_mem\[28\]\[6\] _03934_ _03941_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_184_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_211_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07432_ _02901_ _03075_ _03080_ _02910_ _03081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_51_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_225_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_189_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07363_ _02918_ _02969_ _03012_ _03013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09102_ _04281_ _00713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_31_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06314_ soc.spi_video_ram_1.fifo_in_address\[9\] _02171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_202_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07294_ _02597_ soc.spi_video_ram_1.write_fifo.fifo_mem\[4\]\[10\] _02943_ _02944_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_108_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09033_ _03148_ _04224_ _04240_ _00685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06245_ _02124_ soc.spi_video_ram_1.write_fifo.fifo_mem\[18\]\[2\] _02120_ _02125_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_191_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06176_ soc.rom_encoder_0.sram_sio_oe net53 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_11_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_191_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_172_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09935_ soc.ram_encoder_0.input_bits_left\[2\] _04838_ _04839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_63_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_213_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09866_ soc.cpu.ALU.zx _04741_ _04785_ _04786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_189_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08817_ _03109_ _04124_ _04125_ _00584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_3205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09797_ soc.rom_encoder_0.initializing_step\[3\] _04728_ _04729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_3216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08748_ soc.spi_video_ram_1.write_fifo.fifo_mem\[24\]\[10\] _02411_ _04087_ _04088_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_2515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_199_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1803 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_226_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1814 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1825 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08679_ _04043_ _04046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_81_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1836 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10710_ soc.spi_video_ram_1.fifo_in_address\[6\] _05325_ _05336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_1847 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_42_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1858 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1869 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11690_ _00751_ clknet_leaf_145_wb_clk_i soc.spi_video_ram_1.fifo_in_data\[8\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_214_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_201_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10641_ soc.spi_video_ram_1.write_fifo.fifo_mem\[19\]\[19\] soc.spi_video_ram_1.fifo_in_address\[3\]
+ _05289_ _05299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_41_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10572_ _05256_ _05258_ _01452_ _01207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_6_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12311_ _01339_ clknet_leaf_152_wb_clk_i soc.ram_encoder_0.data_out\[6\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_10_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_177_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_213_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_155_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_170_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12242_ _01270_ clknet_leaf_299_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[29\]\[24\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_5_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_218_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12173_ _01201_ clknet_leaf_126_wb_clk_i soc.boot_loading_offset\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_150_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11124_ _00190_ clknet_leaf_54_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[14\]\[4\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_27_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_231_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_5130 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11055_ _00121_ clknet_leaf_249_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[0\]\[22\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_5141 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5152 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_77_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_236_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5163 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10006_ soc.ram_encoder_0.request_data_out\[6\] soc.ram_encoder_0.data_out\[6\] _04880_
+ _04888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_5174 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5185 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_224_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_218_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3750 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3761 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_229_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3772 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3783 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11957_ _01016_ clknet_leaf_159_wb_clk_i soc.ram_encoder_0.request_data_out\[10\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3794 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_209_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_166_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10908_ soc.spi_video_ram_1.write_fifo.fifo_mem\[8\]\[10\] soc.spi_video_ram_1.fifo_in_data\[10\]
+ _05442_ _05443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_11888_ _00947_ clknet_leaf_318_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[3\]\[14\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_33_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_32_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10839_ _03450_ _05392_ _05405_ _01327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_53_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_158_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_242_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_157_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_203_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06030_ _01908_ _01914_ _01923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_195_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_236_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_177_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_234_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_141_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07981_ soc.spi_video_ram_1.write_fifo.fifo_mem\[0\]\[18\] soc.spi_video_ram_1.write_fifo.fifo_mem\[1\]\[18\]
+ soc.spi_video_ram_1.write_fifo.fifo_mem\[2\]\[18\] soc.spi_video_ram_1.write_fifo.fifo_mem\[3\]\[18\]
+ _02681_ _02758_ _03621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_09720_ _02548_ _02550_ _04685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_101_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_228_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06932_ _02592_ _02593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_41_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_210_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09651_ _04634_ _00910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_28_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06863_ _01717_ _02532_ _02533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_110_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08602_ _04005_ _00489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05814_ _01595_ _01713_ _01714_ soc.cpu.PC.in\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_09582_ _04588_ _04585_ _04589_ _00886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06794_ net66 _02453_ _02472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_243_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08533_ _02122_ soc.spi_video_ram_1.write_fifo.fifo_mem\[2\]\[1\] _03967_ _03969_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_93_1404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_208_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05745_ _01586_ _01649_ _01650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_24_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_169_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_208_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_3_7_0_wb_clk_i clknet_2_3_0_wb_clk_i clknet_3_7_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_24_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08464_ _03930_ _00426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05676_ _01562_ _01583_ _01584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_23_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07415_ soc.spi_video_ram_1.write_fifo.fifo_mem\[14\]\[27\] soc.spi_video_ram_1.write_fifo.fifo_mem\[15\]\[27\]
+ _02613_ _03064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_91_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08395_ _03893_ _00394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_221_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07346_ _02994_ _02995_ _02838_ _02996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_52_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07277_ _02740_ _02927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_163_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09016_ soc.spi_video_ram_1.write_fifo.fifo_mem\[21\]\[18\] _02339_ _04221_ _04232_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_178_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06228_ net62 _02111_ net63 vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_152_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_219_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06159_ _02026_ _02051_ _01454_ _02052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_132_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_1678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09918_ _02111_ _03763_ _04822_ _04825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_28_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_218_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09849_ _04592_ _04761_ _04762_ _04772_ _04773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_98_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_232_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3002 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3013 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_234_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3024 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3035 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_206_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3046 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3057 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xcaravel_hack_soc_97 io_oeb[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_2323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3068 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11811_ _00870_ clknet_leaf_64_wb_clk_i soc.spi_video_ram_1.start_read vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_233_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3079 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_226_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_230_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_183_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11742_ _00803_ clknet_leaf_316_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[4\]\[15\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_183_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11673_ _00734_ clknet_leaf_128_wb_clk_i soc.video_generator_1.v_count\[1\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_39_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_186_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_161_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10624_ _05290_ _01227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_139_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_1395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_6_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10555_ soc.boot_loading_offset\[1\] _05246_ _01395_ _05247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_10_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10486_ soc.cpu.PC.REG.data\[8\] soc.cpu.PC.REG.data\[9\] _05196_ _05203_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_237_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_12225_ _01253_ clknet_leaf_193_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[29\]\[7\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_174_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12156_ _01184_ clknet_leaf_144_wb_clk_i soc.ram_encoder_0.address\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_123_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11107_ _00173_ clknet_leaf_21_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[12\]\[16\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_155_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12087_ soc.cpu.PC.in\[10\] net84 soc.cpu.AReg.data\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_110_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_237_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_211_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_204_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11038_ _00104_ clknet_leaf_226_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[0\]\[5\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_77_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_4270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_225_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_92_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05530_ _01438_ _01440_ _01396_ _00006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_75_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_209_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_36_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2890 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_220_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_178_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07200_ _02849_ _02850_ _02851_ _02852_ _02571_ _02602_ _02853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_08180_ _02165_ soc.spi_video_ram_1.write_fifo.fifo_mem\[10\]\[22\] _03731_ _03756_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_18_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_88_1506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07131_ _02697_ soc.spi_video_ram_1.write_fifo.fifo_mem\[15\]\[4\] _02787_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_118_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_199_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_145_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07062_ _02685_ _02718_ _02720_ _02721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_161_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06013_ _01901_ _01905_ _01906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_12_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_173_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_216_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_141_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_229_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_244_wb_clk_i clknet_5_17_0_wb_clk_i clknet_leaf_244_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_87_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07964_ _02571_ _03604_ _02602_ _03605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_214_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09703_ _04670_ soc.rom_encoder_0.request_address\[12\] _04617_ _04671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_96_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06915_ _00001_ _02576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_114_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_151_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07895_ _02688_ _03537_ _03538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_68_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_216_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09634_ _04625_ _00902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06846_ _02518_ _00221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_83_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_215_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09565_ soc.rom_encoder_0.input_bits_left\[2\] _04575_ _04577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06777_ soc.rom_encoder_0.current_state\[2\] _02435_ _02456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_97_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_93_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_227_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08516_ _02167_ soc.spi_video_ram_1.write_fifo.fifo_mem\[28\]\[23\] _03933_ _03959_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_58_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_212_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05728_ _01595_ _01632_ _01633_ soc.cpu.PC.in\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_09496_ _02250_ soc.cpu.AReg.data\[0\] _04339_ _04533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_149_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_180_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_196_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_169_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08447_ _03921_ _00418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_169_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05659_ _01565_ _01566_ _01567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_211_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_36_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08378_ soc.spi_video_ram_1.write_fifo.fifo_mem\[26\]\[17\] _02337_ _03877_ _03885_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_17_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07329_ _02922_ soc.spi_video_ram_1.write_fifo.fifo_mem\[11\]\[28\] _02722_ _02979_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_178_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_192_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10340_ soc.cpu.ALU.x\[4\] _05109_ _05110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_87_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_191_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10271_ soc.rom_loader.wait_fall_clk soc.rom_loader.writing _05063_ _05064_ _05065_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_105_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12010_ _01069_ clknet_leaf_113_wb_clk_i soc.hack_clock_0.counter\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_191_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_219_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_235_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_207_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2120 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2131 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2142 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2153 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2164 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_199_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2175 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2186 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_202_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11725_ _00786_ clknet_leaf_272_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[9\]\[27\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_leaf_48_wb_clk_i clknet_5_12_0_wb_clk_i clknet_leaf_48_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_1485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_70_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_187_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_175_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11656_ _00717_ clknet_leaf_304_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[20\]\[24\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_70_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_30_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_204_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout90 soc.cpu.AReg.clk net90 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_168_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10607_ _05281_ _01219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_35_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11587_ _00653_ clknet_leaf_241_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[22\]\[23\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_31_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_196_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_182_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10538_ soc.ram_encoder_0.address\[10\] soc.cpu.AReg.data\[10\] _05227_ _05239_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_6_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10469_ soc.cpu.PC.REG.data\[5\] _05186_ _05190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_83_1403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_170_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12208_ _01236_ clknet_leaf_67_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[19\]\[19\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_123_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_233_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_151_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12139_ _01167_ net89 soc.cpu.PC.REG.data\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_97_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_215_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06700_ _02402_ _00191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07680_ _02581_ _03322_ _03325_ _03326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_53_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_168_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_77_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06631_ _02130_ soc.spi_video_ram_1.write_fifo.fifo_mem\[12\]\[5\] _02357_ _02363_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_80_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_94_1532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09350_ soc.rom_encoder_0.write_enable _04426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_06562_ soc.spi_video_ram_1.write_fifo.fifo_mem\[13\]\[5\] _02227_ _02317_ _02323_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_33_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08301_ _03843_ _00350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_61_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_221_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05513_ _01396_ _01427_ _00007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_178_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09281_ _02270_ soc.spi_video_ram_1.write_fifo.fifo_mem\[9\]\[26\] _04359_ _04389_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_181_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06493_ _02128_ soc.spi_video_ram_1.write_fifo.fifo_mem\[0\]\[4\] _02279_ _02284_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_107_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_222_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08232_ _02556_ _03794_ _03795_ _00329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_60_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_159_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08163_ _03747_ _00308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_174_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07114_ soc.spi_video_ram_1.write_fifo.fifo_mem\[24\]\[3\] soc.spi_video_ram_1.write_fifo.fifo_mem\[25\]\[3\]
+ soc.spi_video_ram_1.write_fifo.fifo_mem\[26\]\[3\] soc.spi_video_ram_1.write_fifo.fifo_mem\[27\]\[3\]
+ _02769_ _02770_ _02771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_162_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08094_ _03706_ _00280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_107_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_179_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07045_ _02703_ _02704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_162_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5707 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_134_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5718 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_102_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_5_28_0_wb_clk_i clknet_4_14_0_wb_clk_i clknet_5_28_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XTAP_5729 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08996_ _04220_ _00668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_9_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07947_ _03577_ _03588_ _03579_ _03589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_60_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_217_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07878_ _02656_ _03508_ _03521_ _03522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_244_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09617_ _04612_ _04613_ soc.rom_encoder_0.toggled_sram_sck _04614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_56_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06829_ _02481_ _02485_ _02504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_186_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09548_ _04247_ _04249_ _00878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_184_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_197_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09479_ _04519_ _04522_ _00850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_145_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11510_ _00576_ clknet_leaf_134_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[23\]\[4\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12490_ net49 net48 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_71_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11441_ _00507_ clknet_leaf_269_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[30\]\[22\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_221_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11372_ _00438_ clknet_leaf_36_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[28\]\[11\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_197_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10323_ soc.rom_loader.current_address\[14\] _05098_ _05099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
Xclkbuf_leaf_166_wb_clk_i clknet_5_30_0_wb_clk_i clknet_leaf_166_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_69_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10254_ _03530_ _05044_ _05055_ _01092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_105_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10185_ soc.hack_clock_0.counter\[3\] soc.hack_clock_0.counter\[2\] soc.hack_clock_0.counter\[6\]
+ _05014_ _05015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_121_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_212_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_62_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_234_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_76_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_203_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_230_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_11708_ _00769_ clknet_leaf_17_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[9\]\[10\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_50_1424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11639_ _00700_ clknet_leaf_195_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[20\]\[7\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_50_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xcaravel_hack_soc_190 la_data_out[63] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_237_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08850_ _02311_ _03863_ _04142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_83_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07801_ _02588_ _03442_ _03445_ _03446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_85_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_242_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08781_ _04104_ _00569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_152_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05993_ soc.boot_loading_offset\[1\] _01885_ _01886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_38_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07732_ _03283_ _02625_ _03279_ _03377_ _02734_ _03378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_226_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_211_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07663_ _02902_ _03308_ _03309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_38_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_246_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09402_ soc.rom_encoder_0.output_buffer\[1\] _04460_ _04461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_81_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06614_ _02352_ _00155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_228_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07594_ _02591_ _03240_ _03241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_129_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_244_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_185_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09333_ _04417_ _00808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06545_ _01400_ _01405_ _02311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_179_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_55_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09264_ _04380_ _00776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06476_ soc.spi_video_ram_1.write_fifo.fifo_mem\[16\]\[27\] _02272_ _02216_ _02273_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_08215_ soc.ram_encoder_0.output_buffer\[5\] _02563_ _03783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09195_ soc.spi_video_ram_1.fifo_in_data\[2\] _04341_ _04343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_5_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_146_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08146_ _03738_ _00300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_33_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08077_ soc.spi_video_ram_1.write_fifo.fifo_mem\[11\]\[16\] _02335_ _03691_ _03698_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_134_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07028_ _02685_ _02686_ _02586_ _02687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_6205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_192_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_161_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_216_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_49_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4803 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_130_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4814 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08979_ soc.spi_video_ram_1.write_fifo.fifo_mem\[21\]\[1\] _02393_ _04210_ _04212_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_4825 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4836 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4847 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4858 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11990_ _01049_ clknet_leaf_119_wb_clk_i soc.ram_data_out\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_4869 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10941_ _05459_ _01375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_57_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_216_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10872_ soc.ram_encoder_0.data_out\[10\] _05423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_44_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_232_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_243_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_227_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_242_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_231_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_242_1749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_212_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_164_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_185_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_196_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_123_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11424_ _00490_ clknet_leaf_179_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[30\]\[5\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_184_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_158_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_8 net28 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11355_ _00421_ clknet_leaf_233_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[27\]\[23\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_158_1356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10306_ soc.rom_loader.current_address\[8\] soc.rom_loader.current_address\[7\] _05084_
+ _05088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_98_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11286_ _00352_ clknet_leaf_0_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[1\]\[12\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_79_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_234_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10237_ soc.spi_video_ram_1.fifo_in_data\[13\] _05045_ _05047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_156_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_239_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10168_ soc.ram_encoder_0.initializing_step\[0\] _04919_ soc.ram_encoder_0.initializing_step\[1\]
+ _05002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_120_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10099_ _04846_ _04947_ _04948_ _04949_ _04950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_208_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_212_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_63_wb_clk_i clknet_5_12_0_wb_clk_i clknet_leaf_63_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_235_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_245_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_91_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_231_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06330_ _02113_ soc.spi_video_ram_1.write_fifo.fifo_mem\[17\]\[0\] _02182_ _02183_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_188_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_206_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06261_ _02135_ _00019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_129_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_191_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_141_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08000_ soc.spi_video_ram_1.write_fifo.fifo_mem\[12\]\[17\] soc.spi_video_ram_1.write_fifo.fifo_mem\[13\]\[17\]
+ soc.spi_video_ram_1.write_fifo.fifo_mem\[14\]\[17\] soc.spi_video_ram_1.write_fifo.fifo_mem\[15\]\[17\]
+ _02726_ _03041_ _03639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_102_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06192_ _02077_ _02078_ _02074_ _02079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_191_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_117_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09951_ soc.ram_encoder_0.input_buffer\[1\] _04851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_116_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08902_ soc.spi_video_ram_1.write_fifo.fifo_mem\[25\]\[24\] _04067_ _04143_ _04170_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_135_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09882_ _04609_ _04743_ _04739_ _04797_ _04798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_135_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_217_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08833_ _04133_ _00592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_100_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08764_ soc.spi_video_ram_1.write_fifo.fifo_mem\[24\]\[18\] _02339_ _04087_ _04096_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_3409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05976_ soc.boot_loading_offset\[1\] _01860_ _01862_ _01863_ _01869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_39_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07715_ _02642_ _03353_ _03360_ _02601_ _03361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_39_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2708 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_122_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2719 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08695_ soc.spi_video_ram_1.write_fifo.fifo_mem\[15\]\[17\] _02337_ _04043_ _04057_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_53_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_246_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07646_ _02679_ _03291_ _03292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_57_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_214_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07577_ _02924_ soc.spi_video_ram_1.write_fifo.fifo_mem\[6\]\[13\] _03223_ _02895_
+ _03224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_94_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_41_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_213_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09316_ _02242_ soc.spi_video_ram_1.write_fifo.fifo_mem\[4\]\[12\] _04406_ _04409_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_142_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06528_ _02163_ soc.spi_video_ram_1.write_fifo.fifo_mem\[0\]\[21\] _02278_ _02302_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_224_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_210_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09247_ _04371_ _00768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_107_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_06459_ _02261_ _00091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_222_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_177_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09178_ soc.video_generator_1.v_count\[7\] _04331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_147_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_198_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_159_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08129_ soc.video_generator_1.h_count\[9\] _03727_ _03728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_135_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_190_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11140_ _00206_ clknet_leaf_48_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[14\]\[20\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_1_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_6002 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6013 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput56 net56 io_oeb[24] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_6024 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput67 net67 io_out[19] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_6035 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput78 net78 io_out[35] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_11071_ _00137_ clknet_leaf_202_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[13\]\[9\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_235_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6046 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6057 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6068 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10022_ _04896_ _01019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_6079 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_193_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_5356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_102_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3910 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3921 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3932 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3943 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11973_ _01032_ clknet_leaf_169_wb_clk_i soc.ram_encoder_0.request_address\[10\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_17_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_217_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4699 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3954 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_16_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3965 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3976 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3987 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10924_ soc.spi_video_ram_1.write_fifo.fifo_mem\[8\]\[18\] soc.spi_video_ram_1.fifo_in_address\[2\]
+ _05442_ _05451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_3998 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_186_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10855_ _01613_ _05222_ _05412_ _05414_ _01334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_246_1682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_198_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_213_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10786_ _05376_ _01303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_197_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_207_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_200_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_110_wb_clk_i clknet_5_15_0_wb_clk_i clknet_leaf_110_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_11407_ _00473_ clknet_leaf_78_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[2\]\[17\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_126_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11338_ _00404_ clknet_leaf_201_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[27\]\[6\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_4_9_0_wb_clk_i clknet_3_4_0_wb_clk_i clknet_4_9_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_125_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_154_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11269_ _00335_ clknet_leaf_167_wb_clk_i soc.ram_encoder_0.output_buffer\[15\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_84_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_84_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_39_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_62_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05830_ _01729_ _01730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_23_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5890 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_212_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05761_ _01661_ _01664_ _01585_ _01665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_35_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07500_ soc.spi_video_ram_1.write_fifo.fifo_mem\[21\]\[26\] _03148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_08480_ _03940_ _00432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05692_ soc.ram_data_out\[1\] _01579_ _01599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_169_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07431_ _03076_ _03077_ _03078_ _03079_ _02900_ _03080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_90_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_269_wb_clk_i clknet_5_7_0_wb_clk_i clknet_leaf_269_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_95_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07362_ _02983_ _02992_ _03011_ _02918_ _03012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_52_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09101_ _02258_ soc.spi_video_ram_1.write_fifo.fifo_mem\[20\]\[20\] _04258_ _04281_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06313_ _02170_ _00036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_241_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07293_ _02740_ _02943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_176_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_223_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09032_ _03927_ _04225_ _04240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06244_ soc.spi_video_ram_1.fifo_in_data\[2\] _02124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_190_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_141_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06175_ soc.ram_encoder_0.sram_sio_oe net49 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_137_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09934_ _01378_ _04833_ _04837_ _04838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
X_09865_ _04600_ _04761_ _04762_ _04784_ _04785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_113_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08816_ _04047_ _04124_ _04125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_230_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09796_ soc.rom_encoder_0.initializing_step\[4\] soc.rom_encoder_0.initializing_step\[2\]
+ _04728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_85_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08747_ _04074_ _04087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XTAP_3239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05959_ soc.video_generator_1.v_count\[9\] soc.video_generator_1.v_count\[3\] _01850_
+ _01851_ _01852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or4_1
XTAP_2505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1804 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08678_ _04045_ _00525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_14_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1815 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1826 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_183_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1837 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07629_ _02640_ _03269_ _03275_ _03276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_242_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1859 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10640_ _05298_ _01235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_74_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10571_ soc.hack_wait_clocks\[1\] _05257_ _05258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_122_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_182_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12310_ _01338_ clknet_leaf_154_wb_clk_i soc.ram_encoder_0.data_out\[5\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_195_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12241_ _01269_ clknet_leaf_290_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[29\]\[23\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_202_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_206_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_68_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12172_ _01200_ clknet_leaf_100_wb_clk_i soc.hack_rom_request vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_107_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_194_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_162_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11123_ _00189_ clknet_leaf_54_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[14\]\[3\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_104_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5120 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11054_ _00120_ clknet_leaf_229_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[0\]\[21\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_118_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5131 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_133_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5142 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5153 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10005_ _04887_ _01011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_5164 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5175 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5186 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_5197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3740 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_236_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3751 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3762 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_91_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_209_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_3773 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_opt_4_0_wb_clk_i clknet_5_15_0_wb_clk_i clknet_opt_4_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_11956_ _01015_ clknet_leaf_154_wb_clk_i soc.ram_encoder_0.request_data_out\[9\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3784 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_189_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3795 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10907_ _05429_ _05442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_199_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11887_ _00946_ clknet_leaf_320_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[3\]\[13\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_162_1319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_232_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10838_ soc.spi_video_ram_1.fifo_in_address\[7\] _05393_ _05405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_18_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_186_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10769_ soc.spi_video_ram_1.write_fifo.fifo_mem\[31\]\[20\] soc.spi_video_ram_1.fifo_in_address\[4\]
+ _05355_ _05368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_201_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_186_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_158_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_220_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_113_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07980_ _03577_ _03619_ _03579_ _03620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_99_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_218_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06931_ _02576_ _02592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_84_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_68_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09650_ soc.rom_encoder_0.data_out\[12\] soc.rom_encoder_0.request_data_out\[12\]
+ _04632_ _04634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06862_ _01618_ soc.cpu.AReg.data\[15\] _01718_ soc.ram_data_out\[15\] _02532_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_67_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_228_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08601_ _02128_ soc.spi_video_ram_1.write_fifo.fifo_mem\[30\]\[4\] _04000_ _04005_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_05813_ _01553_ _01669_ soc.cpu.AReg.data\[7\] _01592_ _01714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_110_1410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09581_ net6 _04586_ _04553_ _04589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06793_ soc.rom_encoder_0.output_buffer\[18\] _02455_ _02470_ _02461_ _02471_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_83_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_242_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08532_ _03968_ _00456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_110_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05744_ _01637_ _01646_ _01649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_58_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08463_ soc.spi_video_ram_1.write_fifo.fifo_mem\[27\]\[28\] _02353_ _03898_ _03930_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_224_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05675_ _01563_ _01564_ _01574_ _01582_ soc.cpu.ALU.zy _01583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_1_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_184_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07414_ _03019_ _03040_ _03062_ _03063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_71_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_149_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08394_ soc.spi_video_ram_1.write_fifo.fifo_mem\[26\]\[25\] _02268_ _03865_ _03893_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_52_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07345_ _02703_ soc.spi_video_ram_1.write_fifo.fifo_mem\[16\]\[28\] _02995_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_71_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_192_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_192_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07276_ _02695_ _02926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_192_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_191_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_87_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09015_ _04231_ _00676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06227_ soc.rom_encoder_0.toggled_sram_sck _02111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_121_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06158_ _02027_ _02029_ _02042_ _02050_ _02051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_176_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_160_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_215_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_176_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06089_ soc.video_generator_1.h_count\[1\] soc.video_generator_1.h_count\[2\] _01901_
+ _01982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_236_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09917_ _04821_ _04823_ _04824_ _03714_ _00986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_137_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_246_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_189_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09848_ soc.rom_encoder_0.request_data_out\[7\] _04743_ _04772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_19_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3003 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3014 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3025 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_160_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3036 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_218_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09779_ _04719_ _00953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3047 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3058 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xcaravel_hack_soc_98 io_oeb[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_2324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3069 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11810_ _00010_ clknet_leaf_60_wb_clk_i soc.spi_video_ram_1.fifo_read_request vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11741_ _00802_ clknet_leaf_315_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[4\]\[14\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_214_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_183_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_11672_ _00733_ clknet_leaf_127_wb_clk_i soc.video_generator_1.v_count\[0\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_230_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10623_ soc.spi_video_ram_1.write_fifo.fifo_mem\[19\]\[10\] _02411_ _05289_ _05290_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_161_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_70_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_224_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_183_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10554_ _04243_ _05245_ _05246_ _01201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_155_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10485_ _05171_ _05200_ _05202_ _01175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_170_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_5_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12224_ _01252_ clknet_leaf_211_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[29\]\[6\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_87_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12155_ _01183_ clknet_leaf_144_wb_clk_i soc.ram_encoder_0.address\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_9_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11106_ _00172_ clknet_leaf_3_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[12\]\[15\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_111_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_215_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12086_ soc.cpu.PC.in\[9\] net90 soc.cpu.AReg.data\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_104_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11037_ _00103_ clknet_leaf_200_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[0\]\[4\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_49_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_4260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_224_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_237_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_220_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_166_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_181_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_206_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11939_ _00998_ clknet_leaf_158_wb_clk_i soc.ram_encoder_0.input_buffer\[5\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2880 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2891 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_242_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_222_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_203_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07130_ _02697_ soc.spi_video_ram_1.write_fifo.fifo_mem\[12\]\[4\] _02785_ _02786_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_71_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_179_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_173_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07061_ _02719_ _02720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_103_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06012_ _01902_ _01903_ _01904_ _01905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_161_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_245_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_5_18_0_wb_clk_i clknet_4_9_0_wb_clk_i clknet_5_18_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_88_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07963_ soc.spi_video_ram_1.write_fifo.fifo_mem\[4\]\[19\] soc.spi_video_ram_1.write_fifo.fifo_mem\[5\]\[19\]
+ soc.spi_video_ram_1.write_fifo.fifo_mem\[6\]\[19\] soc.spi_video_ram_1.write_fifo.fifo_mem\[7\]\[19\]
+ _02681_ _02758_ _03604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_9_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_190_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09702_ soc.cpu.PC.REG.data\[12\] soc.rom_loader.current_address\[12\] _04638_ _04670_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06914_ _02574_ _02575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_116_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07894_ soc.spi_video_ram_1.write_fifo.fifo_mem\[9\]\[21\] _03537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_56_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_229_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06845_ soc.rom_encoder_0.output_bits_left\[4\] _02514_ _02517_ _02513_ _02518_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_09633_ soc.rom_encoder_0.data_out\[4\] soc.rom_encoder_0.request_data_out\[4\] _04621_
+ _04625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xclkbuf_leaf_284_wb_clk_i clknet_5_7_0_wb_clk_i clknet_leaf_284_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_167_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_243_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09564_ soc.rom_encoder_0.input_bits_left\[2\] _04575_ _04576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06776_ _02434_ _02454_ _02442_ _02441_ _02455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
Xclkbuf_leaf_213_wb_clk_i clknet_5_20_0_wb_clk_i clknet_leaf_213_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_82_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08515_ _03958_ _00449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05727_ _01553_ soc.cpu.DMuxJMP.sel\[2\] soc.cpu.AReg.data\[2\] _01592_ _01633_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_130_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_230_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09495_ _01387_ _04453_ _01419_ _00856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_208_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08446_ soc.spi_video_ram_1.write_fifo.fifo_mem\[27\]\[20\] _02343_ _03898_ _03921_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_05658_ soc.cpu.AReg.data\[3\] soc.cpu.AReg.data\[2\] _01566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_221_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_212_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_184_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08377_ _03884_ _00385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_177_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05589_ _01488_ _01493_ _01473_ _01497_ _01498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_17_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07328_ _02971_ soc.spi_video_ram_1.write_fifo.fifo_mem\[10\]\[28\] _02978_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_136_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_192_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07259_ _02600_ _02910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_152_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_104_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10270_ soc.rom_encoder_0.write_enable net45 _05064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_118_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_219_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_133_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_239_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_43_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_232_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_246_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_206_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_219_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2110 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2121 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_185_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_15_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_245_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2132 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2143 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_226_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2154 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_167_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2165 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2176 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_1414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2187 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11724_ _00785_ clknet_leaf_281_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[9\]\[26\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11655_ _00716_ clknet_leaf_239_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[20\]\[23\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_243_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10606_ soc.spi_video_ram_1.write_fifo.fifo_mem\[19\]\[2\] _02395_ _05278_ _05281_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_200_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11586_ _00652_ clknet_leaf_240_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[22\]\[22\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_156_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10537_ _05238_ _01192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xclkbuf_leaf_17_wb_clk_i clknet_5_2_0_wb_clk_i clknet_leaf_17_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_171_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10468_ _05171_ _05187_ _05189_ _01171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_174_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12207_ _01235_ clknet_leaf_76_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[19\]\[18\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10399_ _05141_ _01151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_12138_ _01166_ net88 soc.cpu.PC.REG.data\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_229_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_211_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12069_ _01112_ clknet_leaf_111_wb_clk_i soc.rom_loader.current_address\[9\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_78_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_225_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06630_ _02362_ _00161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_4090 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_241_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06561_ _02322_ _00132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_212_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_209_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08300_ _02140_ soc.spi_video_ram_1.write_fifo.fifo_mem\[1\]\[10\] _03842_ _03843_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_05512_ soc.spi_video_ram_1.current_state\[0\] _01397_ _01414_ _01426_ _01427_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_09280_ _03266_ _04375_ _04388_ _00784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06492_ _02283_ _00102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_94_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_146_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08231_ soc.ram_encoder_0.output_buffer\[9\] _02563_ _03795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_147_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08162_ _02147_ soc.spi_video_ram_1.write_fifo.fifo_mem\[10\]\[13\] _03743_ _03747_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_105_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_222_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07113_ _02652_ _02770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_88_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08093_ soc.spi_video_ram_1.write_fifo.fifo_mem\[11\]\[24\] _02266_ _03679_ _03706_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_105_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_134_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_238_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07044_ _02694_ _02703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_133_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_216_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5708 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_88_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5719 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_173_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08995_ soc.spi_video_ram_1.write_fifo.fifo_mem\[21\]\[9\] _02409_ _04210_ _04220_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_29_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07946_ soc.spi_video_ram_1.write_fifo.fifo_mem\[28\]\[20\] soc.spi_video_ram_1.write_fifo.fifo_mem\[29\]\[20\]
+ soc.spi_video_ram_1.write_fifo.fifo_mem\[30\]\[20\] soc.spi_video_ram_1.write_fifo.fifo_mem\[31\]\[20\]
+ _02713_ _02714_ _03588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_151_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07877_ _02640_ _03514_ _03520_ _03521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_151_1395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09616_ soc.hack_rom_request soc.rom_loader.rom_request soc.rom_encoder_0.write_enable
+ _04613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_71_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06828_ soc.ram_encoder_0.output_bits_left\[4\] _02478_ _02503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_83_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_227_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06759_ _02433_ _02437_ _02438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_09547_ _04243_ _04245_ _04246_ _00877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_110_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_231_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_196_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09478_ _01501_ _04521_ _04522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_180_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_211_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_200_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08429_ _03912_ _00409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xclkbuf_4_11_0_wb_clk_i clknet_3_5_0_wb_clk_i clknet_4_11_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_145_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11440_ _00506_ clknet_leaf_231_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[30\]\[21\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_137_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_201_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11371_ _00437_ clknet_leaf_12_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[28\]\[10\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_153_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10322_ soc.rom_loader.current_address\[13\] _05096_ _05098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_180_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10253_ soc.spi_video_ram_1.fifo_in_address\[5\] _05045_ _05055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_1_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_191_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_26_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10184_ _05013_ soc.hack_clock_0.counter\[5\] _05014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_105_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_152_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_135_wb_clk_i clknet_5_24_0_wb_clk_i clknet_leaf_135_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_87_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_212_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_235_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_1506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_207_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_75_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_223_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_15_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_206_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_241_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11707_ _00768_ clknet_leaf_256_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[9\]\[9\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_128_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_163_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_204_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11638_ _00699_ clknet_leaf_210_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[20\]\[6\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_129_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_196_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_171_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11569_ _00635_ clknet_leaf_211_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[22\]\[5\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_6_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_239_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xcaravel_hack_soc_180 la_data_out[53] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_87_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_217_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_171_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xcaravel_hack_soc_191 wbs_ack_o vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_124_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_135_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07800_ _02575_ soc.spi_video_ram_1.write_fifo.fifo_mem\[28\]\[23\] _03444_ _02943_
+ _03445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_170_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08780_ soc.spi_video_ram_1.write_fifo.fifo_mem\[24\]\[26\] _03927_ _04075_ _04104_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_111_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05992_ soc.video_generator_1.v_count\[9\] soc.video_generator_1.v_count\[1\] _01850_
+ _01885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_26_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07731_ _03329_ _03376_ _02918_ _03377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_66_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07662_ soc.spi_video_ram_1.write_fifo.fifo_mem\[9\]\[14\] _03308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_66_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09401_ _04459_ _02460_ _03765_ _02445_ _04460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_65_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06613_ soc.spi_video_ram_1.write_fifo.fifo_mem\[13\]\[27\] _02351_ _02316_ _02352_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_07593_ soc.spi_video_ram_1.write_fifo.fifo_mem\[21\]\[25\] _03240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_213_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09332_ _02258_ soc.spi_video_ram_1.write_fifo.fifo_mem\[4\]\[20\] _04394_ _04417_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06544_ soc.spi_video_ram_1.fifo_in_data\[0\] _02310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_240_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_178_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09263_ _02252_ soc.spi_video_ram_1.write_fifo.fifo_mem\[9\]\[17\] _04359_ _04380_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06475_ soc.spi_video_ram_1.fifo_in_address\[11\] _02272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_166_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08214_ soc.ram_encoder_0.request_address\[4\] _02506_ _03781_ soc.ram_encoder_0.output_buffer\[1\]
+ _03782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_09194_ _00011_ _01613_ _04342_ _00744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_119_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_193_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08145_ _02130_ soc.spi_video_ram_1.write_fifo.fifo_mem\[10\]\[5\] _03732_ _03738_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_135_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08076_ _03697_ _00271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_49_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_162_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07027_ soc.spi_video_ram_1.write_fifo.fifo_mem\[12\]\[2\] soc.spi_video_ram_1.write_fifo.fifo_mem\[13\]\[2\]
+ soc.spi_video_ram_1.write_fifo.fifo_mem\[14\]\[2\] soc.spi_video_ram_1.write_fifo.fifo_mem\[15\]\[2\]
+ _02681_ _02682_ _02686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_6206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_162_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_235_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_130_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_5549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4804 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_118_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4815 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08978_ _04211_ _00659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_4826 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4837 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_217_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4848 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07929_ _02677_ _01392_ _03548_ _03571_ _03572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XTAP_4859 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_244_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10940_ soc.spi_video_ram_1.write_fifo.fifo_mem\[8\]\[26\] _03927_ _05430_ _05459_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_56_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_205_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_186_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_28_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10871_ _01752_ _05221_ _05412_ _05422_ _01342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_72_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_197_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_236_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_223_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_205_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_185_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_5_0_0_wb_clk_i clknet_4_0_0_wb_clk_i clknet_5_0_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_32_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11423_ _00489_ clknet_leaf_197_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[30\]\[4\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_197_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_193_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_9 net34 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11354_ _00420_ clknet_leaf_251_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[27\]\[22\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10305_ soc.rom_loader.current_address\[7\] _05084_ soc.rom_loader.current_address\[8\]
+ _05087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_152_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11285_ _00351_ clknet_leaf_14_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[1\]\[11\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_141_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_316_wb_clk_i clknet_5_0_0_wb_clk_i clknet_leaf_316_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_134_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10236_ _03128_ _05044_ _05046_ _01083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_3_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_171_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10167_ _04999_ _05000_ _05001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_212_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_117_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10098_ soc.ram_encoder_0.request_data_out\[4\] _04930_ _04949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_48_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_222_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_56_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_32_wb_clk_i clknet_5_9_0_wb_clk_i clknet_leaf_32_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_108_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06260_ _02134_ soc.spi_video_ram_1.write_fifo.fifo_mem\[18\]\[7\] _02120_ _02135_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_30_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06191_ _01523_ _01533_ _01528_ _01516_ _02078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_129_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_116_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_171_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09950_ _04846_ _04848_ _04850_ _00993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_08901_ _04169_ _00624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_170_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09881_ soc.rom_encoder_0.request_data_out\[15\] _04742_ _04797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_170_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08832_ _02161_ soc.spi_video_ram_1.write_fifo.fifo_mem\[23\]\[20\] _04109_ _04133_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_98_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05975_ _01852_ _01854_ _01857_ _01867_ _01868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_2
X_08763_ _04095_ _00560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_226_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_211_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07714_ _02581_ _03356_ _03359_ _03360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_38_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_1474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2709 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08694_ _04056_ _00530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_187_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07645_ soc.spi_video_ram_1.write_fifo.fifo_mem\[21\]\[14\] _03291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_53_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07576_ _02907_ _03222_ _03223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_40_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_241_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_55_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09315_ _04408_ _00799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06527_ _02301_ _00119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_22_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06458_ soc.spi_video_ram_1.write_fifo.fifo_mem\[16\]\[21\] _02260_ _02216_ _02261_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_09246_ _02235_ soc.spi_video_ram_1.write_fifo.fifo_mem\[9\]\[9\] _04365_ _04371_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_202_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09177_ _04317_ _04330_ _00739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_215_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06389_ soc.spi_video_ram_1.fifo_in_data\[0\] _02213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_124_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08128_ soc.video_generator_1.h_count\[8\] _03725_ _03727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_107_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08059_ _03688_ _00263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_159_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6003 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput46 net46 io_oeb[10] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_66_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6014 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput57 net57 io_oeb[25] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11070_ _00136_ clknet_leaf_176_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[13\]\[8\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_118_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6025 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput68 net68 io_out[20] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput79 net79 io_out[36] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_6036 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6047 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_6058 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10021_ soc.ram_encoder_0.request_data_out\[13\] soc.ram_encoder_0.data_out\[13\]
+ _04889_ _04896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_66_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6069 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_49_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_88_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3900 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_186_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3911 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3922 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_245_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3933 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11972_ _01031_ clknet_leaf_150_wb_clk_i soc.ram_encoder_0.request_address\[9\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3944 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3955 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3966 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3977 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_1509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10923_ _05450_ _01366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3988 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_147_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3999 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_232_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_204_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10854_ soc.ram_encoder_0.data_out\[1\] _05414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_16_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_227_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_242_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_164_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10785_ soc.spi_video_ram_1.write_fifo.fifo_mem\[31\]\[28\] soc.spi_video_ram_1.fifo_in_address\[12\]
+ _05355_ _05376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_38_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_160_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_125_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11406_ _00472_ clknet_leaf_77_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[2\]\[16\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_201_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11337_ _00403_ clknet_leaf_189_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[27\]\[5\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_leaf_150_wb_clk_i clknet_5_31_0_wb_clk_i clknet_leaf_150_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_98_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_218_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_193_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_158_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_158_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_234_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_175_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11268_ _00334_ clknet_leaf_167_wb_clk_i soc.ram_encoder_0.output_buffer\[14\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_49_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10219_ _05036_ _01076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_11199_ _00265_ clknet_leaf_256_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[11\]\[9\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_121_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_6570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_239_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_228_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5880 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5891 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_208_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05760_ _01662_ _01663_ _01664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_3_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_94_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_235_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05691_ soc.cpu.instruction\[12\] _01598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_36_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_63_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07430_ _02700_ soc.spi_video_ram_1.write_fifo.fifo_mem\[4\]\[27\] _02943_ _03079_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_22_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_223_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_182_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07361_ _02997_ _03003_ _00004_ _03010_ _03011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_91_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_188_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06312_ _02169_ soc.spi_video_ram_1.write_fifo.fifo_mem\[18\]\[24\] _02119_ _02170_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_09100_ _04280_ _00712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_206_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07292_ _02941_ soc.spi_video_ram_1.write_fifo.fifo_mem\[5\]\[10\] _02942_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_104_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09031_ _03240_ _04224_ _04239_ _00684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06243_ _02123_ _00013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_15_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_238_wb_clk_i clknet_5_7_0_wb_clk_i clknet_leaf_238_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_117_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06174_ _02052_ _02066_ _01897_ _01911_ net76 vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_144_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_11_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_190_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09933_ _04834_ _04836_ _04831_ _04837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_176_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_217_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_232_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09864_ soc.rom_encoder_0.request_data_out\[11\] _04742_ _04784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_154_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08815_ _04109_ _04124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_150_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09795_ _04727_ _00961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_73_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_86_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_227_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08746_ _04086_ _00552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05958_ soc.video_generator_1.v_count\[2\] soc.video_generator_1.v_count\[1\] _01851_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XTAP_2506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_213_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05889_ _01705_ _01784_ _01785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08677_ soc.spi_video_ram_1.write_fifo.fifo_mem\[15\]\[11\] _02414_ _04043_ _04045_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_96_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_214_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1816 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1827 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07628_ _02952_ _03272_ _03274_ _03275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_1838 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1849 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07559_ _02707_ _03198_ _03205_ _02970_ _03206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_224_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_210_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10570_ soc.hack_wait_clocks\[0\] _05254_ _05257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_70_1439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_158_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_139_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_194_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09229_ _02219_ soc.spi_video_ram_1.write_fifo.fifo_mem\[9\]\[1\] _04360_ _04362_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_107_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12240_ _01268_ clknet_leaf_269_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[29\]\[22\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_120_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_12171_ _01199_ clknet_leaf_161_wb_clk_i soc.ram_step1_write_request vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_101_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11122_ _00188_ clknet_leaf_54_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[14\]\[2\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_235_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11053_ _00119_ clknet_leaf_51_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[0\]\[20\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_5110 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_172_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5121 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5132 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5143 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10004_ soc.ram_encoder_0.request_data_out\[5\] soc.ram_encoder_0.data_out\[5\] _04880_
+ _04887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_27_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5154 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5165 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5176 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5187 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3730 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_217_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3741 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3752 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3763 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11955_ _01014_ clknet_leaf_154_wb_clk_i soc.ram_encoder_0.request_data_out\[8\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3774 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3785 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_233_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3796 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10906_ _05441_ _01358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_205_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11886_ _00945_ clknet_leaf_1_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[3\]\[12\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_17_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_60_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10837_ _03501_ _05392_ _05404_ _01326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_18_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_207_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10768_ _05367_ _01294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_105_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_200_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10699_ _05330_ _01262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_173_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_218_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_1462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_190_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_68_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_86_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06930_ _02590_ _02591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_113_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_214_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_151_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06861_ _01831_ _02530_ _02531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_83_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08600_ _04004_ _00488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_209_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05812_ _01654_ _01701_ _01712_ _01713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
XFILLER_212_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09580_ soc.rom_encoder_0.input_buffer\[1\] _04588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_06792_ _02443_ _02469_ _02470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_82_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_1591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_188_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_05743_ _01635_ _01647_ _01648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_08531_ _02113_ soc.spi_video_ram_1.write_fifo.fifo_mem\[2\]\[0\] _03967_ _03968_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_149_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_51_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05674_ soc.gpio_i_stored\[0\] _01575_ _01578_ _01581_ _01582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
X_08462_ _03929_ _00425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_23_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07413_ _03046_ _03053_ _03061_ _02655_ _03062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_08393_ _03892_ _00393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_177_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_225_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_189_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07344_ _02712_ soc.spi_video_ram_1.write_fifo.fifo_mem\[17\]\[28\] _02994_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_182_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_143_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_192_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_1286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07275_ _02924_ soc.spi_video_ram_1.write_fifo.fifo_mem\[8\]\[10\] _02925_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_149_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_192_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06226_ _02110_ net73 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09014_ soc.spi_video_ram_1.write_fifo.fifo_mem\[21\]\[17\] _02337_ _04221_ _04231_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_128_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06157_ _02047_ _02049_ _02025_ _02050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_191_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_145_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06088_ _01967_ _01980_ _01924_ _01981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_78_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09916_ soc.rom_encoder_0.initializing_step\[1\] _02459_ soc.rom_encoder_0.initializing_step\[2\]
+ _04824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_24_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_154_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09847_ _04752_ _04771_ _00969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_19_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3004 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_100_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_150_1279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3015 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09778_ _02258_ soc.spi_video_ram_1.write_fifo.fifo_mem\[3\]\[20\] _04696_ _04719_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_3026 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3037 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3048 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3059 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xcaravel_hack_soc_99 io_oeb[8] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_08729_ soc.spi_video_ram_1.write_fifo.fifo_mem\[24\]\[1\] _02393_ _04076_ _04078_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_2336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_215_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11740_ _00801_ clknet_leaf_314_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[4\]\[13\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_242_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11671_ _00732_ clknet_leaf_66_wb_clk_i soc.spi_video_ram_1.state_counter\[10\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10622_ _05276_ _05289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_23_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10553_ _01895_ _05064_ _05246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_6_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_202_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10484_ soc.cpu.PC.in\[9\] _05188_ _05201_ _05202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_108_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12223_ _01251_ clknet_leaf_176_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[29\]\[5\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_154_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_194_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_190_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_174_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12154_ _01182_ clknet_leaf_160_wb_clk_i soc.synch_hack_writeM vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_29_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11105_ _00171_ clknet_leaf_5_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[12\]\[14\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_68_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12085_ soc.cpu.PC.in\[8\] net84 soc.cpu.AReg.data\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_150_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11036_ _00102_ clknet_leaf_199_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[0\]\[3\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_238_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_231_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_213_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_246_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11938_ _00997_ clknet_leaf_158_wb_clk_i soc.ram_encoder_0.input_buffer\[4\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2870 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_127_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2881 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2892 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_232_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11869_ _00928_ clknet_leaf_102_wb_clk_i soc.rom_encoder_0.request_address\[14\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_33_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_193_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_220_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_201_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_158_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_146_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_220_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07060_ _02601_ _02719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_31_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_06011_ soc.video_generator_1.h_count\[2\] _01842_ _01904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_160_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_1249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_142_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07962_ _02768_ _03602_ _03603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09701_ _04669_ _00925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06913_ _02573_ _02574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_64_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07893_ _03021_ soc.spi_video_ram_1.write_fifo.fifo_mem\[11\]\[21\] _02652_ _03536_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_67_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_228_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09632_ _04624_ _00901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06844_ _02445_ _02515_ _02516_ soc.rom_encoder_0.output_bits_left\[4\] _02517_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_95_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09563_ _04565_ _04566_ _04574_ _04575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_110_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06775_ _02433_ _02454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_08514_ _02165_ soc.spi_video_ram_1.write_fifo.fifo_mem\[28\]\[22\] _03933_ _03958_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_05726_ _01615_ _01631_ _01632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_24_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09494_ _02882_ _04532_ _00855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_224_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_184_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08445_ _03920_ _00417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_93_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05657_ soc.cpu.AReg.data\[1\] _01565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_71_1501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_253_wb_clk_i clknet_5_7_0_wb_clk_i clknet_leaf_253_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_145_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_1534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08376_ soc.spi_video_ram_1.write_fifo.fifo_mem\[26\]\[16\] _02335_ _03877_ _03884_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_05588_ _01488_ _01496_ _01497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_108_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_197_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07327_ _02972_ _02973_ _02975_ _02976_ _02642_ _02977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_137_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_197_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07258_ soc.spi_video_ram_1.write_fifo.fifo_mem\[20\]\[9\] soc.spi_video_ram_1.write_fifo.fifo_mem\[21\]\[9\]
+ soc.spi_video_ram_1.write_fifo.fifo_mem\[22\]\[9\] soc.spi_video_ram_1.write_fifo.fifo_mem\[23\]\[9\]
+ _02907_ _02908_ _02909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_136_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06209_ _02092_ _02094_ _02095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_180_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07189_ _02835_ _02837_ _02840_ _02842_ _02656_ _02843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_3_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_28_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_246_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_210_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2100 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2111 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2122 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2133 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2144 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_1726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2155 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2166 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2177 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_243_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_214_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11723_ _00784_ clknet_leaf_239_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[9\]\[25\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_230_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_175_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11654_ _00715_ clknet_leaf_249_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[20\]\[22\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_208_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_202_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10605_ _05280_ _01218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_183_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11585_ _00651_ clknet_leaf_240_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[22\]\[21\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_7_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10536_ soc.ram_encoder_0.address\[9\] soc.cpu.AReg.data\[9\] _05227_ _05238_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_143_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10467_ soc.cpu.PC.in\[5\] _05188_ _05173_ _05189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_155_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_12206_ _01234_ clknet_leaf_79_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[19\]\[17\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_100_1487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10398_ _02248_ soc.spi_video_ram_1.write_fifo.fifo_mem\[6\]\[15\] _05135_ _05141_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_12137_ _01165_ clknet_leaf_163_wb_clk_i soc.cpu.AReg.clk vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_69_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_61_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12068_ _01111_ clknet_leaf_111_wb_clk_i soc.rom_loader.current_address\[8\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_84_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11019_ _00085_ clknet_leaf_10_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[16\]\[15\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_77_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_237_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4080 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4091 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_234_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06560_ soc.spi_video_ram_1.write_fifo.fifo_mem\[13\]\[4\] _02225_ _02317_ _02322_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_94_1534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_206_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05511_ _01418_ _01425_ _01426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06491_ _02126_ soc.spi_video_ram_1.write_fifo.fifo_mem\[0\]\[3\] _02279_ _02283_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_233_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_1589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_205_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_226_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08230_ soc.ram_encoder_0.output_buffer\[5\] _03781_ _03789_ soc.ram_encoder_0.request_data_out\[1\]
+ _03793_ _03794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_127_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08161_ _03746_ _00307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_174_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07112_ _02763_ _02769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_147_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08092_ _03705_ _00279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_140_1278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07043_ _02701_ soc.spi_video_ram_1.write_fifo.fifo_mem\[6\]\[2\] _02702_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_118_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_161_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5709 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_134_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08994_ _04219_ _00667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_64_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07945_ _02678_ _03586_ _03587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_25_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_229_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_214_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07876_ _03515_ _03516_ _03519_ _02723_ _02570_ _03520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_243_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09615_ _02434_ _02447_ _04612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06827_ _02502_ _00218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_55_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09546_ _01396_ _04563_ _00876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06758_ _02434_ _02436_ _02437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_77_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_225_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_221_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05709_ soc.cpu.ALU.no _01615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
X_09477_ _01428_ _04520_ _04521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_164_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06689_ soc.spi_video_ram_1.fifo_in_data\[2\] _02395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_08428_ soc.spi_video_ram_1.write_fifo.fifo_mem\[27\]\[11\] _02414_ _03910_ _03912_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_212_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_205_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08359_ soc.spi_video_ram_1.write_fifo.fifo_mem\[26\]\[8\] _02407_ _03866_ _03875_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_240_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11370_ _00436_ clknet_leaf_256_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[28\]\[9\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_153_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10321_ soc.rom_loader.current_address\[13\] _05096_ _05097_ _01116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_158_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_193_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_69_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10252_ _05054_ _01091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_156_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_65_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_238_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10183_ soc.hack_clock_0.counter\[4\] _05013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_133_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_232_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_219_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_169_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_175_wb_clk_i clknet_5_23_0_wb_clk_i clknet_leaf_175_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_216_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_104_wb_clk_i clknet_5_14_0_wb_clk_i clknet_leaf_104_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_188_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_131_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_215_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_167_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11706_ _00767_ clknet_leaf_178_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[9\]\[8\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_188_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_231_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_188_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_243_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_147_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_198_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11637_ _00698_ clknet_leaf_215_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[20\]\[5\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_180_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11568_ _00634_ clknet_leaf_134_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[22\]\[4\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_171_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10519_ _01564_ _05228_ _05229_ _01183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_143_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11499_ _00565_ clknet_leaf_251_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[24\]\[22\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_87_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_226_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xcaravel_hack_soc_170 la_data_out[43] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xcaravel_hack_soc_181 la_data_out[54] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xcaravel_hack_soc_192 wbs_dat_o[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_130_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_211_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05991_ _01869_ _01872_ _01884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_112_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07730_ _03352_ _03375_ _03376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_22_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_225_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07661_ _02695_ soc.spi_video_ram_1.write_fifo.fifo_mem\[11\]\[14\] _02894_ _03307_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_26_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09400_ _02437_ _02447_ _04459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_1313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_241_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06612_ soc.spi_video_ram_1.fifo_in_address\[11\] _02351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_07592_ _02689_ soc.spi_video_ram_1.write_fifo.fifo_mem\[22\]\[25\] _03238_ _02598_
+ _03239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_207_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_209_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09331_ _04416_ _00807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06543_ _02309_ _00127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_59_1484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09262_ _04379_ _00775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06474_ _02271_ _00096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_244_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08213_ _03780_ _03781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_21_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_194_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_33_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09193_ soc.spi_video_ram_1.fifo_in_data\[1\] _04341_ _04342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_140_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_222_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08144_ _03737_ _00299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_147_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_179_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_140_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08075_ soc.spi_video_ram_1.write_fifo.fifo_mem\[11\]\[15\] _02248_ _03691_ _03697_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_119_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_175_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_235_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07026_ _02596_ _02685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_162_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_162_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_216_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_157_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_118_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_1414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_88_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_130_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_1319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_88_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08977_ soc.spi_video_ram_1.write_fifo.fifo_mem\[21\]\[0\] _02310_ _04210_ _04211_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_195_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4805 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_4816 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4827 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_2_wb_clk_i clknet_5_2_0_wb_clk_i clknet_leaf_2_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_233_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4838 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07928_ _03553_ _03561_ _03570_ _02567_ _03571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_69_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4849 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07859_ _03047_ soc.spi_video_ram_1.write_fifo.fifo_mem\[6\]\[22\] _03502_ _02647_
+ _03503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_56_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10870_ soc.ram_encoder_0.data_out\[9\] _05422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_72_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_244_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_231_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_188_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_164_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09529_ _01451_ _04551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XPHY_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_73_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_200_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_213_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_129_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_184_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_199_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_229_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_201_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11422_ _00488_ clknet_leaf_135_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[30\]\[3\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_126_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_1284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11353_ _00419_ clknet_leaf_233_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[27\]\[21\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_125_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10304_ _05086_ _01110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_10_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11284_ _00350_ clknet_leaf_17_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[1\]\[10\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_112_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10235_ soc.spi_video_ram_1.fifo_in_data\[12\] _05045_ _05046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_80_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10166_ _02548_ _03777_ _05000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_48_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10097_ _04926_ _04948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_130_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_207_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_212_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_223_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_228_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10999_ _00065_ clknet_leaf_301_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[17\]\[24\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_90_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_206_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_241_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_176_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_176_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_1400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06190_ _01471_ _01536_ _01531_ _01519_ _02077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xclkbuf_leaf_72_wb_clk_i clknet_5_9_0_wb_clk_i clknet_leaf_72_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_117_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_239_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_217_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_171_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08900_ soc.spi_video_ram_1.write_fifo.fifo_mem\[25\]\[23\] _04065_ _04143_ _04169_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_09880_ _04787_ _04796_ _00977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_139_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08831_ _04132_ _00591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_98_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08762_ soc.spi_video_ram_1.write_fifo.fifo_mem\[24\]\[17\] _02337_ _04087_ _04095_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_05974_ _01860_ _01866_ _01863_ _01851_ _01867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_66_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07713_ _02783_ soc.spi_video_ram_1.write_fifo.fifo_mem\[4\]\[24\] _03358_ _02741_
+ _03359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_238_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08693_ soc.spi_video_ram_1.write_fifo.fifo_mem\[15\]\[16\] _02335_ _04043_ _04056_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_39_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_199_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07644_ _02703_ soc.spi_video_ram_1.write_fifo.fifo_mem\[23\]\[14\] _02592_ _03290_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_54_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_246_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_226_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_213_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07575_ soc.spi_video_ram_1.write_fifo.fifo_mem\[7\]\[13\] _03222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_81_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09314_ _02240_ soc.spi_video_ram_1.write_fifo.fifo_mem\[4\]\[11\] _04406_ _04408_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_74_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_06526_ _02161_ soc.spi_video_ram_1.write_fifo.fifo_mem\[0\]\[20\] _02278_ _02301_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_90_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_161_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_166_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09245_ _04370_ _00767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06457_ soc.spi_video_ram_1.fifo_in_address\[5\] _02260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_72_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_193_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_182_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_147_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09176_ _01849_ _04328_ _04330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_202_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06388_ _02212_ _00069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_108_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08127_ soc.video_generator_1.h_count\[8\] _03725_ _03726_ _00293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_135_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08058_ soc.spi_video_ram_1.write_fifo.fifo_mem\[11\]\[7\] _02405_ _03680_ _03688_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_66_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6004 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput47 net47 io_oeb[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_150_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07009_ soc.spi_video_ram_1.output_buffer\[22\] _02668_ _02633_ _02669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xoutput58 net58 io_out[10] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_6015 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_6026 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput69 net69 io_out[21] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_6037 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_89_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6048 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10020_ _04895_ _01018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_27_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_231_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6059 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_5336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_118_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_5347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_236_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_76_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3901 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3912 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3923 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11971_ _01030_ clknet_leaf_148_wb_clk_i soc.ram_encoder_0.request_address\[8\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3934 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_56_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_179_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3945 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_205_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_186_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3956 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3967 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10922_ soc.spi_video_ram_1.write_fifo.fifo_mem\[8\]\[17\] soc.spi_video_ram_1.fifo_in_address\[1\]
+ _05442_ _05450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_3978 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3989 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_229_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10853_ _01589_ _05222_ _05412_ _05413_ _01333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_60_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_207_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_201_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10784_ _05375_ _01302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_129_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_185_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_160_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_90_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11405_ _00471_ clknet_leaf_0_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[2\]\[15\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_181_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_236_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11336_ _00402_ clknet_leaf_141_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[27\]\[4\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_154_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11267_ _00333_ clknet_leaf_168_wb_clk_i soc.ram_encoder_0.output_buffer\[13\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_140_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_171_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10218_ _02227_ soc.spi_video_ram_1.write_fifo.fifo_mem\[5\]\[5\] _05030_ _05036_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_6560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11198_ _00264_ clknet_leaf_189_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[11\]\[8\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_122_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_190_wb_clk_i clknet_5_22_0_wb_clk_i clknet_leaf_190_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_6582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10149_ _02484_ _02491_ _02551_ _04987_ _04988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_121_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5870 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_5881 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5892 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_47_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05690_ _01557_ _01596_ _01597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_208_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_184_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_0 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_07360_ _02582_ _03004_ _03009_ _02585_ _03010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_16_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06311_ soc.spi_video_ram_1.fifo_in_address\[8\] _02169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_31_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07291_ _02694_ _02941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_34_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_108_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09030_ _04069_ _04225_ _04239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_30_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_164_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06242_ _02122_ soc.spi_video_ram_1.write_fifo.fifo_mem\[18\]\[1\] _02120_ _02123_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_11_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06173_ _02053_ _02058_ _02059_ _02065_ _02066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_172_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_176_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_117_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_278_wb_clk_i clknet_5_4_0_wb_clk_i clknet_leaf_278_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_132_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09932_ soc.ram_encoder_0.input_bits_left\[2\] _04835_ _04836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_67_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_207_wb_clk_i clknet_5_22_0_wb_clk_i clknet_leaf_207_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_09863_ _04752_ _04783_ _00973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_213_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08814_ _04123_ _00583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_218_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09794_ _02274_ soc.spi_video_ram_1.write_fifo.fifo_mem\[3\]\[28\] _04696_ _04727_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08745_ soc.spi_video_ram_1.write_fifo.fifo_mem\[24\]\[9\] _02409_ _04076_ _04086_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_3219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05957_ soc.video_generator_1.v_count\[8\] soc.video_generator_1.v_count\[7\] _01849_
+ soc.video_generator_1.v_count\[5\] _01850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_4
XFILLER_38_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_242_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_187_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08676_ _04044_ _00524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05888_ _01717_ _01783_ _01784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_26_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1806 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1817 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07627_ _02704_ soc.spi_video_ram_1.write_fifo.fifo_mem\[13\]\[25\] _03273_ _02742_
+ _03274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_1828 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1839 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_241_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_198_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07558_ _02588_ _03201_ _03204_ _03205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_50_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_22_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06509_ _02292_ _00110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_22_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07489_ _02941_ soc.spi_video_ram_1.write_fifo.fifo_mem\[13\]\[12\] _03137_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_202_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09228_ _04361_ _00759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_155_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09159_ soc.video_generator_1.v_count\[0\] _04318_ _04319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_135_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_163_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_237_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12170_ _01198_ clknet_leaf_162_wb_clk_i soc.ram_step2_read_request vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_135_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11121_ _00187_ clknet_leaf_222_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[14\]\[1\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_123_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_122_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_5100 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_7_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11052_ _00118_ clknet_leaf_70_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[0\]\[19\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_5111 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5122 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_5133 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10003_ _04886_ _01010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_7_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5144 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5155 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_237_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5166 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_5177 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3720 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3731 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3742 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3753 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11954_ _01013_ clknet_leaf_153_wb_clk_i soc.ram_encoder_0.request_data_out\[7\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_18_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3764 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3775 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3786 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_232_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3797 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10905_ soc.spi_video_ram_1.write_fifo.fifo_mem\[8\]\[9\] soc.spi_video_ram_1.fifo_in_data\[9\]
+ _05431_ _05441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_166_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11885_ _00944_ clknet_leaf_14_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[3\]\[11\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_242_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10836_ soc.spi_video_ram_1.fifo_in_address\[6\] _05393_ _05404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_220_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10767_ soc.spi_video_ram_1.write_fifo.fifo_mem\[31\]\[19\] soc.spi_video_ram_1.fifo_in_address\[3\]
+ _05355_ _05367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_41_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_146_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_160_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10698_ _02250_ soc.spi_video_ram_1.write_fifo.fifo_mem\[29\]\[16\] _05321_ _05330_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_199_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_201_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_153_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11319_ _00385_ clknet_leaf_19_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[26\]\[16\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12299_ _01327_ clknet_leaf_286_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[7\]\[23\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_leaf_300_wb_clk_i clknet_5_1_0_wb_clk_i clknet_leaf_300_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_49_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_64_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_234_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_171_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_228_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06860_ _01669_ _02529_ _02530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_110_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_110_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05811_ _01669_ _01710_ _01711_ _01712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_227_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06791_ soc.rom_encoder_0.output_buffer\[18\] _02463_ _02464_ soc.rom_encoder_0.request_data_out\[14\]
+ _02469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_23_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08530_ _03966_ _03967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_224_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05742_ _01637_ _01646_ _01647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_36_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08461_ soc.spi_video_ram_1.write_fifo.fifo_mem\[27\]\[27\] _02351_ _03898_ _03929_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_36_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05673_ soc.cpu.instruction\[12\] _01580_ _01581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_223_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07412_ _02901_ _03055_ _03060_ _02910_ _03061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_90_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08392_ soc.spi_video_ram_1.write_fifo.fifo_mem\[26\]\[24\] _02266_ _03865_ _03892_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_149_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07343_ soc.spi_video_ram_1.write_fifo.fifo_mem\[18\]\[28\] soc.spi_video_ram_1.write_fifo.fifo_mem\[19\]\[28\]
+ _02783_ _02993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_71_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_52_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_149_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07274_ _02590_ _02924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_09013_ _04230_ _00675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06225_ _01428_ _01550_ _02110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_145_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06156_ _01921_ _02048_ _02049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_89_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_137_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_06087_ _01925_ _01969_ _01970_ _01980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_104_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_217_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09915_ _02454_ _04731_ _04822_ _04823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_144_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_232_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_154_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09846_ _01615_ _04740_ _04770_ _04771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_63_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_219_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_111_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3005 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_132_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_3016 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09777_ _04718_ _00952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_39_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06989_ _02643_ _02648_ _02649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_3027 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_2_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3038 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3049 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08728_ _04077_ _00543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_214_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08659_ _04035_ _00516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_183_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_199_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_208_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_202_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_183_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11670_ _00731_ clknet_leaf_65_wb_clk_i soc.spi_video_ram_1.state_counter\[9\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_243_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_161_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_224_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_169_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_165_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10621_ _05288_ _01226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_126_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_70_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_183_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_139_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10552_ _04639_ net45 soc.boot_loading_offset\[0\] _05245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_10_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_1349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_211_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10483_ _02053_ _05201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xclkbuf_leaf_129_wb_clk_i clknet_5_12_0_wb_clk_i clknet_leaf_129_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_108_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_185_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12222_ _01250_ clknet_leaf_194_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[29\]\[4\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_13_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_1718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12153_ _01181_ clknet_leaf_162_wb_clk_i soc.hack_clk_strobe vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_68_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_190_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11104_ _00170_ clknet_leaf_16_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[12\]\[13\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_155_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12084_ soc.cpu.PC.in\[7\] net84 soc.cpu.AReg.data\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_2_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11035_ _00101_ clknet_leaf_257_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[0\]\[2\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_77_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_209_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_206_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_233_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11937_ _00996_ clknet_leaf_157_wb_clk_i soc.ram_encoder_0.input_buffer\[3\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_205_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2860 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2871 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2882 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2893 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11868_ _00927_ clknet_5_15_0_wb_clk_i soc.rom_encoder_0.request_address\[13\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_221_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10819_ _03222_ _05392_ _05395_ _01317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_60_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_1484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_207_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11799_ _00859_ clknet_leaf_74_wb_clk_i soc.spi_video_ram_1.fifo_in_address\[2\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_222_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_222_1749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_185_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06010_ soc.video_generator_1.h_count\[1\] _01842_ _01903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_57_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_86_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07961_ soc.spi_video_ram_1.write_fifo.fifo_mem\[0\]\[19\] soc.spi_video_ram_1.write_fifo.fifo_mem\[1\]\[19\]
+ soc.spi_video_ram_1.write_fifo.fifo_mem\[2\]\[19\] soc.spi_video_ram_1.write_fifo.fifo_mem\[3\]\[19\]
+ _02769_ _02770_ _03602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_09700_ _04668_ soc.rom_encoder_0.request_address\[11\] _04617_ _04669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_229_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06912_ _02572_ _02573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_214_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07892_ _02784_ soc.spi_video_ram_1.write_fifo.fifo_mem\[10\]\[21\] _03535_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_68_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09631_ soc.rom_encoder_0.data_out\[3\] soc.rom_encoder_0.request_data_out\[3\] _04621_
+ _04624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_68_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06843_ soc.rom_encoder_0.output_bits_left\[3\] soc.rom_encoder_0.output_bits_left\[2\]
+ _02516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_82_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09562_ _01378_ _04573_ _04574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_3_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06774_ _02438_ _02452_ _02453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_36_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08513_ _03957_ _00448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05725_ _01585_ _01627_ _01630_ _01631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_70_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09493_ soc.spi_video_ram_1.buffer_index\[5\] _04531_ _04532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_36_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08444_ soc.spi_video_ram_1.write_fifo.fifo_mem\[27\]\[19\] _02341_ _03910_ _03920_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_05656_ soc.cpu.AReg.data\[0\] _01564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_2
XFILLER_12_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_225_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_211_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08375_ _03883_ _00384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_56_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05587_ soc.spi_video_ram_1.output_buffer\[1\] _01494_ _01486_ _01495_ _01496_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_162_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07326_ _02577_ _02976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_176_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_293_wb_clk_i clknet_5_4_0_wb_clk_i clknet_leaf_293_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_137_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07257_ _02894_ _02908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_178_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_222_wb_clk_i clknet_5_23_0_wb_clk_i clknet_leaf_222_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_219_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06208_ _02090_ _02093_ _02094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_117_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_238_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07188_ _02643_ _02841_ _02831_ _02842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_121_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_191_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_2_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06139_ _01891_ _01905_ soc.video_generator_1.h_count\[4\] _02031_ _02032_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_133_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_150_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_87_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09829_ soc.rom_encoder_0.request_data_out\[3\] _04743_ _04757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_100_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_150_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2101 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2112 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2123 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_215_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2134 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_161_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2145 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2156 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2167 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_242_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11722_ _00783_ clknet_leaf_276_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[9\]\[24\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_54_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2178 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_203_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11653_ _00714_ clknet_leaf_239_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[20\]\[21\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_74_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_156_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10604_ soc.spi_video_ram_1.write_fifo.fifo_mem\[19\]\[1\] _02393_ _05278_ _05280_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_122_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_204_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11584_ _00650_ clknet_leaf_50_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[22\]\[20\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_126_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_195_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10535_ _05237_ _01191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_13_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_70_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_202_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_109_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10466_ _05170_ _05188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_178_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_12205_ _01233_ clknet_leaf_79_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[19\]\[16\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10397_ _05140_ _01150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xclkbuf_3_6_0_wb_clk_i clknet_2_3_0_wb_clk_i clknet_3_6_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_237_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12136_ _01164_ clknet_leaf_274_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[6\]\[28\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_150_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_215_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_12067_ _01110_ clknet_leaf_111_wb_clk_i soc.rom_loader.current_address\[7\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_leaf_97_wb_clk_i clknet_5_14_0_wb_clk_i clknet_leaf_97_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_133_1242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_238_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11018_ _00084_ clknet_leaf_4_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[16\]\[14\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_77_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_26_wb_clk_i clknet_5_8_0_wb_clk_i clknet_leaf_26_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_168_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4070 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4081 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_4092 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05510_ _01419_ _01423_ _01424_ soc.spi_video_ram_1.current_state\[1\] _01425_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_244_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06490_ _02282_ _00101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_1390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_220_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08160_ _02145_ soc.spi_video_ram_1.write_fifo.fifo_mem\[10\]\[12\] _03743_ _03746_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_105_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07111_ _02767_ _02768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_08091_ soc.spi_video_ram_1.write_fifo.fifo_mem\[11\]\[23\] _02264_ _03679_ _03705_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_147_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07042_ _02700_ _02701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_174_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_173_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_155_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_170_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_192_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08993_ soc.spi_video_ram_1.write_fifo.fifo_mem\[21\]\[8\] _02407_ _04210_ _04219_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_87_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_134_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07944_ soc.spi_video_ram_1.write_fifo.fifo_mem\[24\]\[20\] soc.spi_video_ram_1.write_fifo.fifo_mem\[25\]\[20\]
+ soc.spi_video_ram_1.write_fifo.fifo_mem\[26\]\[20\] soc.spi_video_ram_1.write_fifo.fifo_mem\[27\]\[20\]
+ _02713_ _02714_ _03586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_151_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_68_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_69_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_228_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07875_ _02784_ soc.spi_video_ram_1.write_fifo.fifo_mem\[8\]\[22\] _03518_ _03519_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_29_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_42_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06826_ soc.ram_encoder_0.output_bits_left\[4\] _02495_ _02501_ _02494_ _02502_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_09614_ soc.rom_encoder_0.current_state\[2\] _02457_ _04611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_99_1468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_244_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09545_ soc.spi_video_ram_1.write_fifo.write_pointer\[4\] _04561_ _04563_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_06757_ _02435_ _02436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_71_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_243_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_224_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05708_ _01595_ _01613_ _01614_ soc.cpu.PC.in\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_36_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_58_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09476_ _01379_ soc.spi_video_ram_1.sram_sck_rise_edge _04520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_184_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06688_ _02394_ _00187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_145_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_240_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08427_ _03911_ _00408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_180_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05639_ _01469_ _01542_ _01544_ _01547_ _01548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_24_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08358_ _03874_ _00376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_196_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_7_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07309_ _02954_ _02955_ _02957_ _02958_ _02642_ _02959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_221_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08289_ _02130_ soc.spi_video_ram_1.write_fifo.fifo_mem\[1\]\[5\] _03831_ _03837_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_153_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_203_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10320_ _04426_ soc.rom_loader.was_loading _05096_ soc.rom_loader.current_address\[13\]
+ _05097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_165_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10251_ _02258_ soc.spi_video_ram_1.write_fifo.fifo_mem\[5\]\[20\] _05041_ _05054_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_195_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10182_ soc.hack_clock_0.counter\[0\] _05012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_161_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_94_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_210_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_243_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_128_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_245_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11705_ _00766_ clknet_leaf_191_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[9\]\[7\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_128_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_230_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_144_wb_clk_i clknet_5_28_0_wb_clk_i clknet_leaf_144_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_202_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11636_ _00697_ clknet_leaf_139_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[20\]\[4\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_54_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11567_ _00633_ clknet_leaf_134_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[22\]\[3\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_128_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10518_ soc.ram_encoder_0.address\[0\] _05228_ _05229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_116_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_157_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11498_ _00564_ clknet_leaf_230_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[24\]\[21\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_155_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_171_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xcaravel_hack_soc_160 la_data_out[33] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_100_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_196_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10449_ soc.cpu.PC.REG.data\[0\] soc.cpu.PC.REG.data\[1\] _05175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
Xcaravel_hack_soc_171 la_data_out[44] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xcaravel_hack_soc_182 la_data_out[55] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_152_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xcaravel_hack_soc_193 wbs_dat_o[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_112_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_174_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12119_ _01147_ clknet_leaf_40_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[6\]\[11\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_170_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05990_ _01882_ _01883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_38_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_242_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_187_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07660_ _02783_ soc.spi_video_ram_1.write_fifo.fifo_mem\[10\]\[14\] _03306_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_38_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_226_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_187_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06611_ _02350_ _00154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_81_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07591_ _02591_ _03237_ _03238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_53_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_225_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_46_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_206_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09330_ _02256_ soc.spi_video_ram_1.write_fifo.fifo_mem\[4\]\[19\] _04406_ _04416_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06542_ _02177_ soc.spi_video_ram_1.write_fifo.fifo_mem\[0\]\[28\] _02278_ _02309_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_80_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_222_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_185_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09261_ _02250_ soc.spi_video_ram_1.write_fifo.fifo_mem\[9\]\[16\] _04365_ _04379_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06473_ soc.spi_video_ram_1.write_fifo.fifo_mem\[16\]\[26\] _02270_ _02216_ _02271_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_08212_ _02493_ _03777_ _03779_ _02487_ _03780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_72_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_221_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09192_ _01459_ _04341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_159_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_18_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08143_ _02128_ soc.spi_video_ram_1.write_fifo.fifo_mem\[10\]\[4\] _03732_ _03737_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_119_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08074_ _03696_ _00270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_200_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07025_ _02678_ _02683_ _02684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_150_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_235_1726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08976_ _04209_ _04210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_88_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_4806 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_130_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4817 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_152_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4828 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07927_ _02901_ _03562_ _03569_ _02970_ _03570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_57_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_229_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4839 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07858_ _02700_ _03501_ _03502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_60_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06809_ _02482_ _02485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_16_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07789_ soc.spi_video_ram_1.write_fifo.fifo_mem\[21\]\[23\] _03434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_147_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_225_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09528_ _01430_ _01418_ _01396_ _00871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XPHY_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09459_ _02435_ _04505_ _02524_ _04506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XPHY_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_212_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_90_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_185_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_164_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_240_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_200_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11421_ _00487_ clknet_leaf_261_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[30\]\[2\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_51_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_193_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11352_ _00418_ clknet_leaf_52_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[27\]\[20\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_158_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_193_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_192_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10303_ soc.rom_loader.current_address\[7\] _05084_ _05085_ _05086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_101_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11283_ _00349_ clknet_leaf_248_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[1\]\[9\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_84_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_193_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_238_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10234_ _05029_ _05045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_106_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_161_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10165_ soc.ram_encoder_0.initializing_step\[1\] soc.ram_encoder_0.initializing_step\[0\]
+ _04999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_216_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10096_ _04929_ _04947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_47_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_208_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_169_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_207_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10998_ _00064_ clknet_leaf_233_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[17\]\[23\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_204_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_5_27_0_wb_clk_i clknet_4_13_0_wb_clk_i clknet_5_27_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XTAP_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_143_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_231_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_188_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_30_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_203_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11619_ _00685_ clknet_leaf_287_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[21\]\[26\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_50_1246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_204_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_190_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_1448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_1702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_67_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_41_wb_clk_i clknet_5_6_0_wb_clk_i clknet_leaf_41_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_174_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08830_ _02159_ soc.spi_video_ram_1.write_fifo.fifo_mem\[23\]\[19\] _04109_ _04132_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_97_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08761_ _04094_ _00559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05973_ soc.video_generator_1.v_count\[0\] _01866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XTAP_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_230_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07712_ _02679_ _03357_ _03358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08692_ _03404_ _04046_ _04055_ _00529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_54_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_96_1405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07643_ _02893_ soc.spi_video_ram_1.write_fifo.fifo_mem\[22\]\[14\] _03289_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_96_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_183_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_207_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07574_ soc.spi_video_ram_1.write_fifo.fifo_mem\[0\]\[13\] soc.spi_video_ram_1.write_fifo.fifo_mem\[1\]\[13\]
+ soc.spi_video_ram_1.write_fifo.fifo_mem\[2\]\[13\] soc.spi_video_ram_1.write_fifo.fifo_mem\[3\]\[13\]
+ _03139_ _02895_ _03221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_59_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_41_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09313_ _04407_ _00798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_94_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06525_ _02300_ _00118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_161_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_22_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_228_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09244_ _02233_ soc.spi_video_ram_1.write_fifo.fifo_mem\[9\]\[8\] _04365_ _04370_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_146_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06456_ _02259_ _00090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_142_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09175_ _04317_ _04329_ _00738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_222_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06387_ _02177_ soc.spi_video_ram_1.write_fifo.fifo_mem\[17\]\[28\] _02181_ _02212_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_08126_ _01959_ _03712_ _03725_ soc.video_generator_1.h_count\[8\] _01380_ _03726_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_179_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_174_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08057_ _03687_ _00262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_116_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07008_ _02627_ _02667_ _02668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_6005 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput48 net48 io_oeb[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_162_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_153_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6016 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput59 net59 io_out[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_6027 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_88_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6038 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6049 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_5326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_89_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_5337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_131_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_5348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_233_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_188_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08959_ soc.spi_video_ram_1.write_fifo.fifo_mem\[22\]\[21\] _04061_ _04177_ _04201_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_4636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3902 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_4658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3913 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3924 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11970_ _01029_ clknet_leaf_147_wb_clk_i soc.ram_encoder_0.request_address\[7\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_91_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3935 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3946 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3957 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10921_ _05449_ _01365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_245_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3968 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_147_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3979 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_244_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10852_ soc.ram_encoder_0.data_out\[0\] _05413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_186_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_73_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_241_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_188_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10783_ soc.spi_video_ram_1.write_fifo.fifo_mem\[31\]\[27\] soc.spi_video_ram_1.fifo_in_address\[11\]
+ _05355_ _05375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XPHY_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_213_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_184_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_199_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_201_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_201_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11404_ _00470_ clknet_leaf_320_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[2\]\[14\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_138_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11335_ _00401_ clknet_leaf_140_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[27\]\[3\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_99_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11266_ _00332_ clknet_leaf_168_wb_clk_i soc.ram_encoder_0.output_buffer\[12\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_45_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10217_ _05035_ _01075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_136_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11197_ _00263_ clknet_leaf_192_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[11\]\[7\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_6561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_234_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10148_ _02548_ _04917_ _04987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_6594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5860 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_5871 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_23_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5882 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5893 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10079_ soc.ram_data_out\[0\] _04927_ _04933_ _04934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_78_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_212_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_236_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_1 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_225_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_211_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_206_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_147_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_1534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_225_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06310_ _02168_ _00035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_108_1545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07290_ _02744_ soc.spi_video_ram_1.write_fifo.fifo_mem\[6\]\[10\] _02895_ _02940_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_87_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06241_ soc.spi_video_ram_1.fifo_in_data\[1\] _02122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_223_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_191_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06172_ _01903_ _02060_ _02063_ _02064_ _02065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_102_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09931_ soc.ram_encoder_0.input_bits_left\[3\] soc.ram_encoder_0.input_bits_left\[4\]
+ _04835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_144_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_154_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09862_ _01702_ _04741_ _04782_ _04783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08813_ _02143_ soc.spi_video_ram_1.write_fifo.fifo_mem\[23\]\[11\] _04117_ _04123_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_246_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09793_ _04726_ _00960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_189_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_247_wb_clk_i clknet_5_19_0_wb_clk_i clknet_leaf_247_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_85_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_3209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08744_ _04085_ _00551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05956_ soc.video_generator_1.v_count\[6\] _01849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_27_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08675_ soc.spi_video_ram_1.write_fifo.fifo_mem\[15\]\[10\] _02411_ _04043_ _04044_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_2519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_199_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05887_ _01618_ soc.cpu.AReg.data\[12\] _01718_ soc.ram_data_out\[12\] _01783_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_22_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_226_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_183_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1807 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07626_ _02931_ soc.spi_video_ram_1.write_fifo.fifo_mem\[12\]\[25\] _03273_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_1818 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1829 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_242_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07557_ _02924_ soc.spi_video_ram_1.write_fifo.fifo_mem\[28\]\[13\] _03203_ _02927_
+ _03204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_201_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06508_ _02143_ soc.spi_video_ram_1.write_fifo.fifo_mem\[0\]\[11\] _02290_ _02292_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_166_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07488_ soc.spi_video_ram_1.write_fifo.fifo_mem\[8\]\[12\] soc.spi_video_ram_1.write_fifo.fifo_mem\[9\]\[12\]
+ soc.spi_video_ram_1.write_fifo.fifo_mem\[10\]\[12\] soc.spi_video_ram_1.write_fifo.fifo_mem\[11\]\[12\]
+ _02574_ _02577_ _03136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_50_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06439_ soc.spi_video_ram_1.fifo_in_data\[15\] _02248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_09227_ _02213_ soc.spi_video_ram_1.write_fifo.fifo_mem\[9\]\[0\] _04360_ _04361_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_182_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_6_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09158_ _01959_ _03712_ _04318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_107_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_194_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_202_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08109_ _03714_ _01968_ _03715_ _00286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_135_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09089_ _02246_ soc.spi_video_ram_1.write_fifo.fifo_mem\[20\]\[14\] _04270_ _04275_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_11_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_218_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11120_ _00186_ clknet_leaf_178_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[14\]\[0\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_66_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11051_ _00117_ clknet_leaf_76_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[0\]\[18\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_66_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_231_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5101 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5112 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5123 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10002_ soc.ram_encoder_0.request_data_out\[4\] soc.ram_encoder_0.data_out\[4\] _04880_
+ _04886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_118_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5134 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5145 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_191_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_190_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_77_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_236_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5156 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5167 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5178 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3710 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3721 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_4477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3732 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3743 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_218_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11953_ _01012_ clknet_leaf_152_wb_clk_i soc.ram_encoder_0.request_data_out\[6\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3754 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3765 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3776 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_229_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3787 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10904_ _05440_ _01357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3798 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11884_ _00943_ clknet_leaf_17_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[3\]\[10\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_60_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_207_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10835_ _03527_ _05392_ _05403_ _01325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_246_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_158_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_53_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10766_ _05366_ _01293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_242_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_186_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10697_ _03396_ _05324_ _05329_ _01261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_160_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11318_ _00384_ clknet_leaf_314_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[26\]\[15\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_113_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_12298_ _01326_ clknet_leaf_268_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[7\]\[22\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_141_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11249_ _00315_ clknet_leaf_52_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[10\]\[20\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_64_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_41_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_68_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_6391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05810_ _01704_ _01709_ _01711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_67_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06790_ _02453_ _02467_ _02468_ _01381_ _00215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_5690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05741_ _01562_ _01645_ _01646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_242_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_208_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_1408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08460_ _03928_ _00424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_58_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05672_ soc.ram_data_out\[0\] _01579_ _01580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07411_ _02578_ _03057_ _03058_ _03059_ _02900_ _03060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_224_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08391_ _03891_ _00392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_56_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_177_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07342_ _02655_ _02991_ _02992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_148_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_221_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07273_ _02922_ soc.spi_video_ram_1.write_fifo.fifo_mem\[11\]\[10\] _02647_ _02923_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_164_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09012_ soc.spi_video_ram_1.write_fifo.fifo_mem\[21\]\[16\] _02335_ _04221_ _04230_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_136_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06224_ _02096_ _02107_ _02109_ _01428_ net72 vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_163_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_195_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_145_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06155_ _01922_ _02004_ _02048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_176_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_219_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06086_ _01924_ _01978_ _01979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09914_ soc.rom_encoder_0.initializing_step\[2\] soc.rom_encoder_0.initializing_step\[1\]
+ _02459_ _04822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_154_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09845_ _04590_ _04761_ _04762_ _04769_ _04770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_115_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_218_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3006 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09776_ _02256_ soc.spi_video_ram_1.write_fifo.fifo_mem\[3\]\[19\] _04708_ _04718_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_39_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06988_ soc.spi_video_ram_1.write_fifo.fifo_mem\[0\]\[1\] soc.spi_video_ram_1.write_fifo.fifo_mem\[1\]\[1\]
+ soc.spi_video_ram_1.write_fifo.fifo_mem\[2\]\[1\] soc.spi_video_ram_1.write_fifo.fifo_mem\[3\]\[1\]
+ _02645_ _02647_ _02648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_3017 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3028 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_160_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3039 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08727_ soc.spi_video_ram_1.write_fifo.fifo_mem\[24\]\[0\] _02310_ _04076_ _04077_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_05939_ _01682_ _01827_ _01831_ _01832_ _01833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_27_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08658_ soc.spi_video_ram_1.write_fifo.fifo_mem\[15\]\[2\] _02395_ _04032_ _04035_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_226_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_4_8_0_wb_clk_i clknet_3_4_0_wb_clk_i clknet_4_8_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XTAP_1626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_241_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_230_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07609_ soc.spi_video_ram_1.write_fifo.fifo_mem\[5\]\[25\] _03256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_42_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_169_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_148_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_168_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08589_ _03997_ _00484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_168_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10620_ soc.spi_video_ram_1.write_fifo.fifo_mem\[19\]\[9\] _02409_ _05278_ _05288_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_41_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_243_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10551_ _05063_ _05244_ _01200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_183_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10482_ soc.cpu.PC.REG.data\[9\] _05199_ _05200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_155_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12221_ _01249_ clknet_leaf_139_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[29\]\[3\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_204_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_237_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12152_ _01180_ net89 soc.cpu.PC.REG.data\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_174_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_1749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_169_wb_clk_i clknet_5_31_0_wb_clk_i clknet_leaf_169_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_151_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11103_ _00169_ clknet_leaf_7_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[12\]\[12\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12083_ soc.cpu.PC.in\[6\] net84 soc.cpu.AReg.data\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_133_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11034_ _00100_ clknet_leaf_215_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[0\]\[1\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_89_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_237_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_49_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_77_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_224_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11936_ _00995_ clknet_leaf_160_wb_clk_i soc.ram_encoder_0.input_buffer\[2\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2850 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2861 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_206_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_166_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2872 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_127_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2883 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11867_ _00926_ clknet_leaf_104_wb_clk_i soc.rom_encoder_0.request_address\[12\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2894 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_220_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10818_ soc.spi_video_ram_1.fifo_in_data\[13\] _05393_ _05395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_186_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11798_ _00858_ clknet_leaf_83_wb_clk_i soc.spi_video_ram_1.fifo_in_address\[1\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_41_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_203_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_146_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10749_ soc.spi_video_ram_1.write_fifo.fifo_mem\[31\]\[11\] soc.spi_video_ram_1.fifo_in_data\[11\]
+ _05355_ _05357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_118_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_199_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_177_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_141_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07960_ _03577_ _03600_ _03579_ _03601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_99_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06911_ _00000_ _02572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_136_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07891_ _02767_ _03526_ _03533_ _02910_ _03534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_151_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09630_ _04623_ _00900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_99_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06842_ _02434_ _02435_ _02515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_28_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09561_ _04567_ _04571_ soc.rom_encoder_0.toggled_sram_sck _04572_ _04573_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_06773_ _02448_ _02451_ _02452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_23_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_243_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05724_ _01585_ _01629_ _01630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08512_ _02163_ soc.spi_video_ram_1.write_fifo.fifo_mem\[28\]\[21\] _03933_ _03957_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_110_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09492_ _01460_ _01464_ _04520_ _04524_ _04531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_227_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_223_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_212_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05655_ soc.cpu.instruction\[12\] _01563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_149_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08443_ _03919_ _00416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_196_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08374_ soc.spi_video_ram_1.write_fifo.fifo_mem\[26\]\[15\] _02248_ _03877_ _03883_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_149_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05586_ soc.spi_video_ram_1.output_buffer\[3\] soc.spi_video_ram_1.output_buffer\[2\]
+ _01461_ _01495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_143_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_20_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07325_ _02696_ soc.spi_video_ram_1.write_fifo.fifo_mem\[12\]\[28\] _02974_ _02975_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_71_1558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07256_ _02679_ _02907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_197_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_192_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06207_ _01470_ _01485_ _01463_ _02093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07187_ soc.spi_video_ram_1.write_fifo.fifo_mem\[8\]\[6\] soc.spi_video_ram_1.write_fifo.fifo_mem\[9\]\[6\]
+ soc.spi_video_ram_1.write_fifo.fifo_mem\[10\]\[6\] soc.spi_video_ram_1.write_fifo.fifo_mem\[11\]\[6\]
+ _02680_ _02722_ _02841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
Xclkbuf_opt_3_0_wb_clk_i clknet_5_15_0_wb_clk_i clknet_opt_3_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_238_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06138_ soc.video_generator_1.h_count\[7\] _02031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_132_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_156_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xclkbuf_leaf_262_wb_clk_i clknet_5_7_0_wb_clk_i clknet_leaf_262_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_191_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06069_ _01945_ _01958_ _01960_ _01962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_59_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_232_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_235_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_219_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09828_ _04752_ _04756_ _00965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_86_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_246_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_235_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_206_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_189_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09759_ _04709_ _00943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2102 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2113 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2124 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2135 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2146 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2157 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_167_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2168 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_199_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_1406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11721_ _00782_ clknet_leaf_238_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[9\]\[23\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2179 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_202_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11652_ _00713_ clknet_leaf_51_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[20\]\[20\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_23_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10603_ _05279_ _01217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_128_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11583_ _00649_ clknet_leaf_29_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[22\]\[19\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10534_ soc.ram_encoder_0.address\[8\] soc.cpu.AReg.data\[8\] _05227_ _05237_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_10_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_156_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_196_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10465_ soc.cpu.PC.REG.data\[5\] _05186_ _05187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_6_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12204_ _01232_ clknet_leaf_10_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[19\]\[15\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10396_ _02246_ soc.spi_video_ram_1.write_fifo.fifo_mem\[6\]\[14\] _05135_ _05140_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_151_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12135_ _01163_ clknet_leaf_273_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[6\]\[27\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_123_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_111_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12066_ _01109_ clknet_leaf_108_wb_clk_i soc.rom_loader.current_address\[6\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_137_1390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_81_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11017_ _00083_ clknet_leaf_11_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[16\]\[13\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_65_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4060 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_225_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4071 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4082 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4093 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_66_wb_clk_i clknet_5_11_0_wb_clk_i clknet_leaf_66_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_205_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11919_ _00978_ clknet_leaf_121_wb_clk_i soc.cpu.instruction\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_33_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_221_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1990 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_207_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_222_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_140_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07110_ _02706_ _02767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_53_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08090_ _03704_ _00278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_101_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07041_ _02644_ _02700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_122_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_1722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08992_ _04218_ _00666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_115_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_233_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_229_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07943_ _03576_ _03580_ _03582_ _03584_ _02710_ _03585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_214_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_155_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_205_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07874_ _02712_ _03517_ _03518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_217_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09613_ _04609_ _04586_ _04610_ _00896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_84_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06825_ soc.ram_encoder_0.output_bits_left\[4\] _02496_ _02497_ _02500_ _02501_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_3_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09544_ _04562_ _00875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_06756_ soc.rom_encoder_0.current_state\[1\] _02435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_70_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05707_ _01553_ soc.cpu.DMuxJMP.sel\[1\] soc.cpu.AReg.data\[1\] _01592_ _01614_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_06687_ soc.spi_video_ram_1.write_fifo.fifo_mem\[14\]\[1\] _02393_ _02391_ _02394_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_09475_ _02674_ _04517_ _04518_ _01392_ _04519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_34_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_24_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_197_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08426_ soc.spi_video_ram_1.write_fifo.fifo_mem\[27\]\[10\] _02411_ _03910_ _03911_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_05638_ _01519_ _01545_ _01546_ _01471_ soc.spi_video_ram_1.buffer_index\[4\] _01547_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_211_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_200_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_162_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05569_ _01468_ soc.spi_video_ram_1.output_buffer\[12\] _01477_ soc.spi_video_ram_1.output_buffer\[13\]
+ _01478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_08357_ soc.spi_video_ram_1.write_fifo.fifo_mem\[26\]\[7\] _02405_ _03866_ _03874_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_165_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07308_ _02577_ _02958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_123_1467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08288_ _03836_ _00344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_109_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_197_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07239_ soc.spi_video_ram_1.write_fifo.fifo_mem\[4\]\[9\] soc.spi_video_ram_1.write_fifo.fifo_mem\[5\]\[9\]
+ soc.spi_video_ram_1.write_fifo.fifo_mem\[6\]\[9\] soc.spi_video_ram_1.write_fifo.fifo_mem\[7\]\[9\]
+ _02712_ _02722_ _02890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_125_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_238_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10250_ _05053_ _01090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_152_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10181_ soc.ram_encoder_0.initializing_step\[4\] _05010_ _05011_ _01063_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_117_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_212_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_207_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_234_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_203_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_5_17_0_wb_clk_i clknet_4_8_0_wb_clk_i clknet_5_17_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XTAP_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11704_ _00765_ clknet_leaf_205_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[9\]\[6\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_187_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11635_ _00696_ clknet_leaf_139_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[20\]\[3\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_129_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_204_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11566_ _00632_ clknet_leaf_55_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[22\]\[2\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_leaf_184_wb_clk_i clknet_5_29_0_wb_clk_i clknet_leaf_184_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_156_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_183_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10517_ _05227_ _05228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_11497_ _00563_ clknet_leaf_261_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[24\]\[20\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_109_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_113_wb_clk_i clknet_5_26_0_wb_clk_i clknet_leaf_113_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_87_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xcaravel_hack_soc_150 la_data_out[22] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_10448_ soc.cpu.PC.REG.data\[0\] _05171_ _05174_ _01166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xcaravel_hack_soc_161 la_data_out[34] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xcaravel_hack_soc_172 la_data_out[45] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_124_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xcaravel_hack_soc_183 la_data_out[56] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_237_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xcaravel_hack_soc_194 wbs_dat_o[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_112_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10379_ _02229_ soc.spi_video_ram_1.write_fifo.fifo_mem\[6\]\[6\] _05124_ _05131_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_124_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12118_ _01146_ clknet_leaf_15_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[6\]\[10\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_97_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_215_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_238_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12049_ net26 clknet_leaf_173_wb_clk_i soc.rom_encoder_0.data_out\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_38_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06610_ soc.spi_video_ram_1.write_fifo.fifo_mem\[13\]\[26\] _02270_ _02316_ _02350_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_07590_ soc.spi_video_ram_1.write_fifo.fifo_mem\[23\]\[25\] _03237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_52_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_168_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_228_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06541_ _02308_ _00126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_94_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_244_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06472_ soc.spi_video_ram_1.fifo_in_address\[10\] _02270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_09260_ _03410_ _04375_ _04378_ _00774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_181_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08211_ _03778_ _03779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09191_ _04340_ _00743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_147_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08142_ _03736_ _00298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_179_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08073_ soc.spi_video_ram_1.write_fifo.fifo_mem\[11\]\[14\] _02246_ _03691_ _03696_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_140_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_140_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07024_ soc.spi_video_ram_1.write_fifo.fifo_mem\[8\]\[2\] soc.spi_video_ram_1.write_fifo.fifo_mem\[9\]\[2\]
+ soc.spi_video_ram_1.write_fifo.fifo_mem\[10\]\[2\] soc.spi_video_ram_1.write_fifo.fifo_mem\[11\]\[2\]
+ _02681_ _02682_ _02683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_128_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_162_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_192_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_5519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08975_ _02311_ _04175_ _04209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_9_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_60_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4807 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4818 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07926_ _02642_ _03565_ _03568_ _03569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_4829 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_151_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07857_ soc.spi_video_ram_1.write_fifo.fifo_mem\[7\]\[22\] _03501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_17_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_244_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_216_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06808_ soc.ram_encoder_0.current_state\[2\] _02484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_28_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_147_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07788_ _02689_ soc.spi_video_ram_1.write_fifo.fifo_mem\[22\]\[23\] _03432_ _02598_
+ _03433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_71_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09527_ _02673_ _04549_ _04550_ _03714_ _00870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_06739_ _02425_ _00207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_77_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_240_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_73_1439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09458_ soc.rom_encoder_0.request_data_out\[9\] _02441_ _04505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_227_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_08409_ soc.spi_video_ram_1.write_fifo.fifo_mem\[27\]\[2\] _02395_ _03899_ _03902_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_12_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09389_ soc.spi_video_ram_1.state_sram_clk_counter\[2\] soc.spi_video_ram_1.state_sram_clk_counter\[1\]
+ soc.spi_video_ram_1.state_sram_clk_counter\[3\] _04452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_196_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_205_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11420_ _00486_ clknet_leaf_222_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[30\]\[1\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_138_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11351_ _00417_ clknet_leaf_35_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[27\]\[19\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_117_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10302_ soc.rom_loader.current_address\[7\] _05084_ _05070_ _05085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_3_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11282_ _00348_ clknet_leaf_220_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[1\]\[8\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_84_1535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10233_ _05041_ _05044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_161_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_234_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10164_ _04998_ _01058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10095_ _04787_ _04946_ _01041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_43_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_235_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_90_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10997_ _00063_ clknet_leaf_267_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[17\]\[22\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_245_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_108_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_230_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11618_ _00684_ clknet_leaf_241_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[21\]\[25\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_54_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11549_ _00615_ clknet_leaf_318_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[25\]\[14\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_176_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_144_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_143_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_174_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_170_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_4_10_0_wb_clk_i clknet_3_5_0_wb_clk_i clknet_4_10_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_112_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_135_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_239_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08760_ soc.spi_video_ram_1.write_fifo.fifo_mem\[24\]\[16\] _02335_ _04087_ _04094_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_112_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05972_ _01859_ _01864_ _01865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_81_wb_clk_i clknet_5_10_0_wb_clk_i clknet_leaf_81_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_113_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07711_ soc.spi_video_ram_1.write_fifo.fifo_mem\[5\]\[24\] _03357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_66_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08691_ _04054_ _04048_ _04055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_66_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_226_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_211_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xclkbuf_leaf_10_wb_clk_i clknet_5_3_0_wb_clk_i clknet_leaf_10_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_93_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_1488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07642_ _02958_ _03284_ _03287_ _02706_ _03288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_96_1439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07573_ _02831_ _03213_ _03219_ _03220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_41_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_222_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_185_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09312_ _02237_ soc.spi_video_ram_1.write_fifo.fifo_mem\[4\]\[10\] _04406_ _04407_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06524_ _02159_ soc.spi_video_ram_1.write_fifo.fifo_mem\[0\]\[19\] _02290_ _02300_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_94_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09243_ _04369_ _00766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06455_ soc.spi_video_ram_1.write_fifo.fifo_mem\[16\]\[20\] _02258_ _02216_ _02259_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_221_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_210_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06386_ _02211_ _00068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09174_ _01939_ _04326_ _04328_ _04329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_194_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_1426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08125_ _03713_ _03724_ _03725_ _00292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_198_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_200_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08056_ soc.spi_video_ram_1.write_fifo.fifo_mem\[11\]\[6\] _02403_ _03680_ _03687_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_190_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07007_ _02606_ _02657_ _02666_ _02667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_6006 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_157_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput49 net49 io_oeb[13] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_6017 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_118_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_6028 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_235_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6039 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_49_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_130_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08958_ _04200_ _00650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_4615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_69_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_243_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_229_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3903 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07909_ _03550_ _03551_ _02976_ _03552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_44_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3914 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3925 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08889_ _04163_ _00618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_5_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_245_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_3936 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3947 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10920_ soc.spi_video_ram_1.write_fifo.fifo_mem\[8\]\[16\] soc.spi_video_ram_1.fifo_in_address\[0\]
+ _05442_ _05449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_217_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3958 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_16_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3969 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_245_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_246_1620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_246_1631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10851_ _05411_ _05412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_38_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_72_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_198_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10782_ _03157_ _05358_ _05374_ _01301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_242_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_212_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_164_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_234_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_197_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_240_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_200_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11403_ _00469_ clknet_leaf_319_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[2\]\[13\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_184_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_177_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11334_ _00400_ clknet_leaf_195_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[27\]\[2\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_177_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_141_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_238_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11265_ _00331_ clknet_leaf_169_wb_clk_i soc.ram_encoder_0.output_buffer\[11\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_158_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_180_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_1313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10216_ _02225_ soc.spi_video_ram_1.write_fifo.fifo_mem\[5\]\[4\] _05030_ _05035_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_80_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11196_ _00262_ clknet_leaf_203_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[11\]\[6\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_6551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10147_ _04873_ _04925_ _04986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_94_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5850 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5861 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5872 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_11_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_1753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5883 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10078_ _04928_ _04931_ _04932_ _04933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_94_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_5894 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_208_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_95_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_204_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_91_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_231_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_188_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_203_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06240_ _02121_ _00012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_54_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06171_ _01949_ _01947_ _01959_ _01842_ _02064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_190_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09930_ _02480_ _02498_ _04834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_172_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09861_ _04598_ _04761_ _04762_ _04781_ _04782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08812_ _04122_ _00582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_112_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_154_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09792_ _02272_ soc.spi_video_ram_1.write_fifo.fifo_mem\[3\]\[27\] _04696_ _04726_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_230_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08743_ soc.spi_video_ram_1.write_fifo.fifo_mem\[24\]\[8\] _02407_ _04076_ _04085_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_05955_ _01841_ _01847_ _01848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_41_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_227_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_213_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08674_ _04031_ _04043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_96_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05886_ _01702_ _01781_ _01782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_66_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_287_wb_clk_i clknet_5_5_0_wb_clk_i clknet_leaf_287_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_57_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07625_ _03047_ soc.spi_video_ram_1.write_fifo.fifo_mem\[14\]\[25\] _03271_ _02593_
+ _03272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_1808 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1819 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_183_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_216_wb_clk_i clknet_5_21_0_wb_clk_i clknet_leaf_216_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_41_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07556_ _02907_ _03202_ _03203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_59_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_228_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06507_ _02291_ _00109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07487_ _02984_ _03127_ _03134_ _02601_ _03135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_42_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_179_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_206_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09226_ _04359_ _04360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_107_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_241_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06438_ _02247_ _00084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_72_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09157_ _01939_ _02034_ _04316_ _01380_ _04317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_4
XFILLER_33_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06369_ _02159_ soc.spi_video_ram_1.write_fifo.fifo_mem\[17\]\[19\] _02193_ _02203_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_159_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08108_ _01926_ _01994_ _03715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_135_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09088_ _04274_ _00706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08039_ _03596_ _03675_ _03676_ _00255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_107_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_194_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_239_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11050_ _00116_ clknet_leaf_78_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[0\]\[17\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_153_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5102 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5113 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_89_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10001_ _04885_ _01009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_103_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5124 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_133_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5135 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5146 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5157 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5168 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5179 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_184_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_4445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3700 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3711 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3722 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3733 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11952_ _01011_ clknet_leaf_153_wb_clk_i soc.ram_encoder_0.request_data_out\[5\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3744 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3755 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_45_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3766 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3777 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10903_ soc.spi_video_ram_1.write_fifo.fifo_mem\[8\]\[8\] soc.spi_video_ram_1.fifo_in_data\[8\]
+ _05431_ _05440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_244_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3788 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3799 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11883_ _00942_ clknet_leaf_249_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[3\]\[9\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_83_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_246_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_199_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10834_ soc.spi_video_ram_1.fifo_in_address\[5\] _05393_ _05403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_57_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_246_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_232_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_213_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10765_ soc.spi_video_ram_1.write_fifo.fifo_mem\[31\]\[18\] soc.spi_video_ram_1.fifo_in_address\[2\]
+ _05355_ _05366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_40_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_199_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_186_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_201_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10696_ soc.spi_video_ram_1.fifo_in_data\[15\] _05325_ _05329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_51_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_172_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_185_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_220_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11317_ _00383_ clknet_leaf_318_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[26\]\[14\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_126_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12297_ _01325_ clknet_leaf_292_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[7\]\[21\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_107_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11248_ _00314_ clknet_leaf_30_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[10\]\[19\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_136_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_45_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_218_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11179_ _00245_ clknet_leaf_60_wb_clk_i soc.spi_video_ram_1.output_buffer\[11\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_6381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_110_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_23_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_209_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_212_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_1583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05740_ _01598_ soc.cpu.AReg.data\[3\] _01639_ _01644_ _01606_ _01645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_236_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4990 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_149_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05671_ soc.cpu.AReg.data\[14\] soc.cpu.AReg.data\[13\] _01579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_36_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07410_ _02700_ soc.spi_video_ram_1.write_fifo.fifo_mem\[6\]\[11\] _02577_ _03059_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_23_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08390_ soc.spi_video_ram_1.write_fifo.fifo_mem\[26\]\[23\] _02264_ _03865_ _03891_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_91_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_189_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_182_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07341_ _02984_ _02985_ _02990_ _02601_ _02991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_149_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07272_ _02695_ _02922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_192_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_223_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_192_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09011_ _03387_ _04224_ _04229_ _00674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_148_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06223_ _01485_ _01475_ _02108_ _02109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_191_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06154_ _01978_ _02045_ _02046_ _02047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_89_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06085_ _01972_ _01974_ _01977_ _01978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_144_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09913_ soc.rom_encoder_0.initializing_step\[2\] _04818_ _04821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_236_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_160_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09844_ soc.rom_encoder_0.request_data_out\[6\] _04743_ _04769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_58_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_74_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09775_ _04717_ _00951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06987_ _02646_ _02647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_3007 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3018 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_6_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08726_ _04075_ _04076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XTAP_3029 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05938_ _01682_ _01822_ _01825_ _01832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_2306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_226_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08657_ _04034_ _00515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_163_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05869_ _01654_ _01766_ _01767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_81_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07608_ soc.spi_video_ram_1.write_fifo.fifo_mem\[0\]\[25\] soc.spi_video_ram_1.write_fifo.fifo_mem\[1\]\[25\]
+ soc.spi_video_ram_1.write_fifo.fifo_mem\[2\]\[25\] soc.spi_video_ram_1.write_fifo.fifo_mem\[3\]\[25\]
+ _02680_ _02838_ _03255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_42_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_242_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_187_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08588_ _02177_ soc.spi_video_ram_1.write_fifo.fifo_mem\[2\]\[28\] _03966_ _03997_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_42_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_214_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07539_ soc.spi_video_ram_1.output_buffer\[11\] _02676_ _03187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_10_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10550_ _05218_ soc.hack_clk_strobe _05244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_224_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09209_ _00011_ _01736_ _04350_ _00751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_154_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10481_ soc.cpu.PC.REG.data\[8\] _05196_ _05199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_167_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12220_ _01248_ clknet_leaf_262_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[29\]\[2\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_202_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_191_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12151_ _01179_ net89 soc.cpu.PC.REG.data\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_136_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_151_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11102_ _00168_ clknet_leaf_38_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[12\]\[11\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_215_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12082_ soc.cpu.PC.in\[5\] net89 soc.cpu.AReg.data\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_81_1313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11033_ _00099_ clknet_leaf_219_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[0\]\[0\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_215_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_leaf_138_wb_clk_i clknet_5_25_0_wb_clk_i clknet_leaf_138_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_213_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_218_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11935_ _00994_ clknet_leaf_158_wb_clk_i soc.ram_encoder_0.input_buffer\[1\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_27_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_245_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2840 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_79_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2851 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2862 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2873 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11866_ _00925_ clknet_leaf_104_wb_clk_i soc.rom_encoder_0.request_address\[11\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_60_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2884 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_177_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2895 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10817_ _03131_ _05392_ _05394_ _01316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_14_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11797_ _00857_ clknet_leaf_82_wb_clk_i soc.spi_video_ram_1.fifo_in_address\[0\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_14_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_242_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10748_ _05356_ _01285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_179_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10679_ _02233_ soc.spi_video_ram_1.write_fifo.fifo_mem\[29\]\[8\] _05310_ _05319_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_160_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_154_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12349_ _01377_ clknet_leaf_278_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[8\]\[28\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_47_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06910_ _02570_ _02571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_9_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07890_ _02582_ _03529_ _03532_ _03533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_60_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_190_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06841_ soc.rom_encoder_0.output_bits_left\[3\] _02513_ _02514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_67_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09560_ soc.rom_encoder_0.request_write _02462_ _04565_ _04572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_7_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06772_ _02437_ _02450_ _02451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_83_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_237_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08511_ _03956_ _00447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_110_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_208_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05723_ _01617_ _01626_ _01628_ _01629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_184_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09491_ _01460_ _04520_ _04530_ _04519_ _00854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_36_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08442_ soc.spi_video_ram_1.write_fifo.fifo_mem\[27\]\[18\] _02339_ _03910_ _03919_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_110_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_224_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_208_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05654_ _01561_ _01562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_91_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08373_ _03882_ _00383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05585_ _01461_ soc.spi_video_ram_1.buffer_index\[1\] _01494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_108_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_221_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07324_ _02590_ soc.spi_video_ram_1.write_fifo.fifo_mem\[13\]\[28\] _02974_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_104_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_220_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_197_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_143_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07255_ _02901_ _02905_ _02906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_149_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_165_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06206_ _01487_ _01490_ _01491_ _01486_ _02087_ _02092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_121_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07186_ _02570_ _02839_ _02840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_180_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06137_ _01930_ _01931_ _01940_ _02030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_133_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_219_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06068_ _01945_ _01958_ _01960_ _01961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_87_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09827_ soc.cpu.DMuxJMP.sel\[2\] _04740_ _04755_ _04756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_232_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_leaf_231_wb_clk_i clknet_5_5_0_wb_clk_i clknet_leaf_231_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_228_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09758_ _02237_ soc.spi_video_ram_1.write_fifo.fifo_mem\[3\]\[10\] _04708_ _04709_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_246_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2103 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08709_ soc.spi_video_ram_1.fifo_in_address\[7\] _04065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_2114 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2125 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_227_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09689_ _04660_ soc.rom_encoder_0.request_address\[8\] _04617_ _04661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_2136 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2147 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2158 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11720_ _00781_ clknet_leaf_238_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[9\]\[22\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_230_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2169 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_243_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_163_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11651_ _00712_ clknet_leaf_32_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[20\]\[19\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10602_ soc.spi_video_ram_1.write_fifo.fifo_mem\[19\]\[0\] soc.spi_video_ram_1.fifo_in_data\[0\]
+ _05278_ _05279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_11_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_243_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11582_ _00648_ clknet_leaf_27_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[22\]\[18\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_196_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout84 net85 net84 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_141_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_183_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_161_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10533_ _05236_ _01190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_7_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_210_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_155_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10464_ soc.cpu.PC.REG.data\[4\] _05183_ _05186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_183_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_237_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_12203_ _01231_ clknet_leaf_3_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[19\]\[14\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_164_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10395_ _05139_ _01149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_48_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12134_ _01162_ clknet_leaf_295_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[6\]\[26\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_97_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_319_wb_clk_i clknet_5_0_0_wb_clk_i clknet_leaf_319_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_61_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_12065_ _01108_ clknet_leaf_112_wb_clk_i soc.rom_loader.current_address\[5\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_237_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11016_ _00082_ clknet_leaf_4_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[16\]\[12\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_211_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4050 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4061 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4072 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_219_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4083 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4094 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_185_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_206_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11918_ _00977_ clknet_leaf_121_wb_clk_i soc.cpu.instruction\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_18_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_209_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_220_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2692 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_127_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11849_ _00908_ clknet_leaf_87_wb_clk_i soc.rom_encoder_0.request_data_out\[10\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_53_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1980 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1991 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_202_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_35_wb_clk_i clknet_5_9_0_wb_clk_i clknet_leaf_35_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_105_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_70_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07040_ _02697_ soc.spi_video_ram_1.write_fifo.fifo_mem\[5\]\[2\] _02698_ _02699_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_62_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_161_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_216_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08991_ soc.spi_video_ram_1.write_fifo.fifo_mem\[21\]\[7\] _02405_ _04210_ _04218_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_138_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07942_ _02571_ _03583_ _02602_ _03584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_60_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07873_ soc.spi_video_ram_1.write_fifo.fifo_mem\[9\]\[22\] _03517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_84_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_233_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09612_ soc.rom_encoder_0.input_buffer\[7\] _04584_ _04601_ _04610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_110_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06824_ _02498_ _02499_ _02500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_68_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_243_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09543_ _04254_ _04560_ _04561_ _04562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_209_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06755_ soc.rom_encoder_0.current_state\[2\] _02434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_4
XFILLER_83_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_227_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05706_ _01556_ _01612_ _01613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_221_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_212_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09474_ _01378_ _01410_ _04518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_225_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06686_ soc.spi_video_ram_1.fifo_in_data\[1\] _02393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_164_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_196_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08425_ _03897_ _03910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_05637_ soc.spi_video_ram_1.output_buffer\[6\] soc.spi_video_ram_1.output_buffer\[7\]
+ _01467_ _01546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_36_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08356_ _03873_ _00375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05568_ _01461_ _01476_ _01477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_165_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07307_ _02941_ soc.spi_video_ram_1.write_fifo.fifo_mem\[20\]\[10\] _02956_ _02957_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_138_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08287_ _02128_ soc.spi_video_ram_1.write_fifo.fifo_mem\[1\]\[4\] _03831_ _03836_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_192_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05499_ soc.spi_video_ram_1.start_read _01408_ _01412_ _01413_ _01414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_166_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07238_ _02643_ _02888_ _02889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_124_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07169_ soc.spi_video_ram_1.write_fifo.fifo_mem\[16\]\[6\] soc.spi_video_ram_1.write_fifo.fifo_mem\[17\]\[6\]
+ soc.spi_video_ram_1.write_fifo.fifo_mem\[18\]\[6\] soc.spi_video_ram_1.write_fifo.fifo_mem\[19\]\[6\]
+ _02645_ _02614_ _02823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_30_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_191_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10180_ _02482_ _05003_ _05010_ soc.ram_encoder_0.initializing_step\[4\] _01380_
+ _05011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_65_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_238_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_121_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_219_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_235_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_199_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_131_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_231_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_202_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_188_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11703_ _00764_ clknet_leaf_222_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[9\]\[5\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_54_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11634_ _00695_ clknet_leaf_137_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[20\]\[2\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_141_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11565_ _00631_ clknet_leaf_208_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[22\]\[1\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_10_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_196_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10516_ _05226_ _05227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_116_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11496_ _00562_ clknet_leaf_34_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[24\]\[19\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_143_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xcaravel_hack_soc_140 la_data_out[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_10447_ soc.cpu.PC.in\[0\] _05172_ _05173_ _05174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xcaravel_hack_soc_151 la_data_out[23] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_152_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xcaravel_hack_soc_162 la_data_out[35] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_87_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xcaravel_hack_soc_173 la_data_out[46] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_170_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xcaravel_hack_soc_184 la_data_out[57] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_83_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_217_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xcaravel_hack_soc_195 wbs_dat_o[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_10378_ _05130_ _01141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_112_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_153_wb_clk_i clknet_5_30_0_wb_clk_i clknet_leaf_153_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_2_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12117_ _01145_ clknet_leaf_249_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[6\]\[9\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_112_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12048_ net25 clknet_opt_1_0_wb_clk_i soc.rom_encoder_0.data_out\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_26_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_238_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_225_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_187_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_81_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_19_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06540_ _02175_ soc.spi_video_ram_1.write_fifo.fifo_mem\[0\]\[27\] _02278_ _02308_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_3190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_207_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_228_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_221_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06471_ _02269_ _00095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_34_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08210_ _02484_ _02491_ _02479_ _03778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_60_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_222_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09190_ _02213_ _04338_ _04339_ _04340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_92_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_187_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_147_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08141_ _02126_ soc.spi_video_ram_1.write_fifo.fifo_mem\[10\]\[3\] _03732_ _03736_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_18_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08072_ _03695_ _00269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_31_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_162_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_179_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07023_ _02598_ _02682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_235_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_157_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08974_ _04208_ _00658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_29_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4808 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07925_ _02635_ soc.spi_video_ram_1.write_fifo.fifo_mem\[30\]\[21\] _03567_ _02904_
+ _03568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_60_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4819 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_217_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07856_ soc.spi_video_ram_1.write_fifo.fifo_mem\[0\]\[22\] soc.spi_video_ram_1.write_fifo.fifo_mem\[1\]\[22\]
+ soc.spi_video_ram_1.write_fifo.fifo_mem\[2\]\[22\] soc.spi_video_ram_1.write_fifo.fifo_mem\[3\]\[22\]
+ _02700_ _02647_ _03500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_112_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06807_ _02480_ _02481_ _02482_ _02483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_186_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07787_ _02591_ _03431_ _03432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_44_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09526_ soc.spi_video_ram_1.start_read _02673_ _04550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06738_ soc.spi_video_ram_1.write_fifo.fifo_mem\[14\]\[21\] _02260_ _02390_ _02425_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_213_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_73_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_197_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09457_ _02445_ _02441_ _04459_ _04504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XPHY_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_06669_ _02382_ _00180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_52_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_200_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_08408_ _03901_ _00399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_129_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09388_ _04451_ _00829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_244_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08339_ soc.spi_video_ram_1.write_fifo.write_pointer\[4\] _01403_ _03862_ _03863_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_138_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11350_ _00416_ clknet_leaf_23_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[27\]\[18\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_197_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10301_ _05071_ _05083_ _05084_ _01109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_153_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_180_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_158_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11281_ _00347_ clknet_leaf_205_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[1\]\[7\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_4_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10232_ _05043_ _01082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_105_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10163_ _04831_ _04993_ _04994_ _02484_ _01395_ _04998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_0_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_82_1282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_212_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10094_ soc.ram_data_out\[3\] _04927_ _04945_ _04946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_87_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_134_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_207_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_112_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_21_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_1722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10996_ _00062_ clknet_leaf_235_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[17\]\[21\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_128_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_203_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_241_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_187_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_176_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_223_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_204_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_145_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11617_ _00683_ clknet_leaf_303_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[21\]\[24\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_156_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_102_1327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11548_ _00614_ clknet_leaf_315_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[25\]\[13\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_183_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_184_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_239_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11479_ _00545_ clknet_leaf_196_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[24\]\[2\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_171_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_05971_ _01860_ _01861_ _01862_ _01863_ _01864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_25_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07710_ _02783_ soc.spi_video_ram_1.write_fifo.fifo_mem\[6\]\[24\] _03355_ _02894_
+ _03356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_66_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08690_ soc.spi_video_ram_1.fifo_in_data\[15\] _04054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_07641_ _03285_ _03286_ _02690_ _03287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_187_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_246_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_228_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07572_ _02582_ _03216_ _03218_ _03219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_50_wb_clk_i clknet_5_6_0_wb_clk_i clknet_leaf_50_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_62_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09311_ _04393_ _04406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_22_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06523_ _02299_ _00117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_179_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09242_ _02231_ soc.spi_video_ram_1.write_fifo.fifo_mem\[9\]\[7\] _04365_ _04369_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06454_ soc.spi_video_ram_1.fifo_in_address\[4\] _02258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_241_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09173_ _01939_ _02034_ _04325_ _04328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_06385_ _02175_ soc.spi_video_ram_1.write_fifo.fifo_mem\[17\]\[27\] _02181_ _02211_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_202_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08124_ soc.video_generator_1.h_count\[7\] _03723_ _03725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_147_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_124_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_194_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_162_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08055_ _03686_ _00261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_134_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07006_ _02659_ _02661_ _02663_ _02665_ _02620_ _02666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_89_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_192_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_190_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6007 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6018 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6029 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_143_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_5317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08957_ soc.spi_video_ram_1.write_fifo.fifo_mem\[22\]\[20\] _02343_ _04177_ _04200_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_88_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07908_ _02926_ soc.spi_video_ram_1.write_fifo.fifo_mem\[16\]\[21\] _03551_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_4649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3904 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08888_ soc.spi_video_ram_1.write_fifo.fifo_mem\[25\]\[17\] _02337_ _04155_ _04163_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_3915 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3926 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_244_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3937 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3948 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07839_ _02607_ _03482_ _03483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_99_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3959 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10850_ _05219_ _05244_ _05411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_232_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_246_1643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09509_ _04539_ _00863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_10781_ _03927_ _05359_ _05374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_227_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_201_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_158_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_73_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_160_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_205_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_227_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11402_ _00468_ clknet_leaf_1_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[2\]\[12\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_165_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11333_ _00399_ clknet_leaf_188_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[27\]\[1\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_181_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_153_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11264_ _00330_ clknet_leaf_169_wb_clk_i soc.ram_encoder_0.output_buffer\[10\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_218_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_234_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10215_ _05034_ _01074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_49_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_2_3_0_wb_clk_i clknet_0_wb_clk_i clknet_2_3_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XTAP_6530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_171_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11195_ _00261_ clknet_leaf_207_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[11\]\[5\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_6541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_95_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_239_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10146_ _03714_ _04985_ _01053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_6574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5840 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_79_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_5851 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_5862 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_236_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5873 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10077_ net1 _04834_ _04932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_5884 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5895 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_235_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_169_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_3 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_44_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_245_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10979_ _00045_ clknet_leaf_140_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[17\]\[4\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_225_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_182_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_54_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06170_ _02061_ _01902_ _01903_ _02062_ _02063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_184_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_158_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_193_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09860_ soc.rom_encoder_0.request_data_out\[10\] _04742_ _04781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_63_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_217_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08811_ _02140_ soc.spi_video_ram_1.write_fifo.fifo_mem\[23\]\[10\] _04117_ _04122_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_113_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09791_ _04725_ _00959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08742_ _04084_ _00550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05954_ _01844_ _01846_ _01847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_61_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_226_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08673_ _04042_ _00523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05885_ _01670_ soc.cpu.ALU.x\[12\] _01781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_113_1286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07624_ _02613_ _03270_ _03271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_214_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07555_ soc.spi_video_ram_1.write_fifo.fifo_mem\[29\]\[13\] _03202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_81_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_241_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06506_ _02140_ soc.spi_video_ram_1.write_fifo.fifo_mem\[0\]\[10\] _02290_ _02291_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_224_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07486_ _02706_ _03130_ _03133_ _03134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_39_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_210_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_256_wb_clk_i clknet_5_18_0_wb_clk_i clknet_leaf_256_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_09225_ _04358_ _04359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_06437_ soc.spi_video_ram_1.write_fifo.fifo_mem\[16\]\[14\] _02246_ _02238_ _02247_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_194_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09156_ soc.video_generator_1.v_count\[2\] _04314_ _04315_ _04316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_147_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06368_ _02202_ _00059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_198_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08107_ _01395_ _03714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_09087_ _02244_ soc.spi_video_ram_1.write_fifo.fifo_mem\[20\]\[13\] _04270_ _04274_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_163_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06299_ soc.spi_video_ram_1.fifo_in_address\[4\] _02161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_163_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_163_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08038_ soc.spi_video_ram_1.output_buffer\[1\] _02675_ _03676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_190_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_235_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5103 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10000_ soc.ram_encoder_0.request_data_out\[3\] soc.ram_encoder_0.data_out\[3\] _04880_
+ _04885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_153_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5114 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_172_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5125 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_130_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5136 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_114_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09989_ _02504_ _04873_ _04877_ _04878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XTAP_4402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_114_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5147 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5158 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_218_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5169 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_44_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3701 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3712 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3723 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11951_ _01010_ clknet_leaf_155_wb_clk_i soc.ram_encoder_0.request_data_out\[4\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3734 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_217_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3745 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3756 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3767 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10902_ _05439_ _01356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3778 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11882_ _00941_ clknet_leaf_216_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[3\]\[8\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_233_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3789 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10833_ _05402_ _01324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_198_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_242_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10764_ _05365_ _01292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_164_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_197_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_200_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10695_ _03300_ _05324_ _05328_ _01260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_55_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_201_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_103_1488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11316_ _00382_ clknet_leaf_315_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[26\]\[13\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12296_ _01324_ clknet_leaf_49_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[7\]\[20\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_180_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11247_ _00313_ clknet_leaf_25_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[10\]\[18\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_190_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11178_ _00244_ clknet_leaf_60_wb_clk_i soc.spi_video_ram_1.output_buffer\[12\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_94_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_171_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10129_ soc.ram_data_out\[11\] _04928_ _04972_ _04973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_5670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_95_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_208_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5692 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4980 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4991 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05670_ net77 _01564_ _01576_ _01577_ _01578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_169_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_223_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07340_ _02986_ _02987_ _02988_ _02989_ _02900_ _02990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_188_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_225_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07271_ _02920_ soc.spi_video_ram_1.write_fifo.fifo_mem\[10\]\[10\] _02921_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09010_ _04054_ _04225_ _04229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06222_ soc.spi_video_ram_1.buffer_index\[4\] _02090_ soc.spi_video_ram_1.buffer_index\[5\]
+ _02108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_129_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06153_ _01924_ _02046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_145_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_172_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06084_ _01976_ _01906_ _01977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_172_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09912_ _04817_ _04820_ _00985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_176_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_232_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09843_ _04752_ _04768_ _00968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_99_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_150_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_230_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06986_ _02576_ _02646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09774_ _02254_ soc.spi_video_ram_1.write_fifo.fifo_mem\[3\]\[18\] _04708_ _04717_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_80_1583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3008 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3019 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_227_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05937_ _01828_ _01829_ _01830_ _01831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_08725_ _04074_ _04075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_167_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08656_ soc.spi_video_ram_1.write_fifo.fifo_mem\[15\]\[1\] _02393_ _04032_ _04034_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_05868_ _01682_ _01763_ _01764_ _01765_ _01766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_82_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_215_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_167_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_183_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_148_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07607_ _03236_ _03244_ _03253_ _02567_ _03254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_82_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_208_1722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08587_ _03996_ _00483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05799_ _01595_ _01699_ _01700_ soc.cpu.PC.in\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_109_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_228_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_1411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_243_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07538_ _01419_ _03107_ _03185_ _02677_ _03186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_165_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_179_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07469_ soc.spi_video_ram_1.write_fifo.fifo_mem\[24\]\[12\] soc.spi_video_ram_1.write_fifo.fifo_mem\[25\]\[12\]
+ soc.spi_video_ram_1.write_fifo.fifo_mem\[26\]\[12\] soc.spi_video_ram_1.write_fifo.fifo_mem\[27\]\[12\]
+ _03054_ _02904_ _03117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_122_1319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09208_ soc.spi_video_ram_1.fifo_in_data\[8\] _04346_ _04350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_10480_ _05171_ _05197_ _05198_ _01174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_120_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09139_ soc.spi_video_ram_1.state_counter\[6\] _04302_ _04304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_108_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_136_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12150_ _01178_ net89 soc.cpu.PC.REG.data\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_194_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11101_ _00167_ clknet_leaf_16_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[12\]\[10\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_78_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12081_ soc.cpu.PC.in\[4\] net84 soc.cpu.AReg.data\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_151_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11032_ _00098_ clknet_leaf_277_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[16\]\[28\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_77_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_76_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_77_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11934_ _00993_ clknet_leaf_158_wb_clk_i soc.ram_encoder_0.input_buffer\[0\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2830 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2841 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2852 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_178_wb_clk_i clknet_5_23_0_wb_clk_i clknet_leaf_178_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_3597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_205_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2863 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11865_ _00924_ clknet_leaf_109_wb_clk_i soc.rom_encoder_0.request_address\[10\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2874 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2885 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2896 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_232_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_107_wb_clk_i clknet_5_15_0_wb_clk_i clknet_leaf_107_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_10816_ soc.spi_video_ram_1.fifo_in_data\[12\] _05393_ _05394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_18_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11796_ _00856_ clknet_leaf_71_wb_clk_i soc.spi_video_ram_1.sram_sio_oe vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_43_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10747_ soc.spi_video_ram_1.write_fifo.fifo_mem\[31\]\[10\] soc.spi_video_ram_1.fifo_in_data\[10\]
+ _05355_ _05356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_201_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_159_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_12_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10678_ _05318_ _01253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_185_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_220_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_51_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12348_ _01376_ clknet_leaf_271_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[8\]\[27\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_173_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_181_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12279_ _01307_ clknet_leaf_262_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[7\]\[3\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_68_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_218_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06840_ _01379_ _02456_ _02448_ _02513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_110_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_231_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_209_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06771_ _02433_ _02449_ _02450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_83_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_236_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08510_ _02161_ soc.spi_video_ram_1.write_fifo.fifo_mem\[28\]\[20\] _03933_ _03956_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_05722_ _01560_ _01584_ _01609_ _01608_ _01597_ _01628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_2
XFILLER_48_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_97_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09490_ _01428_ _01465_ _04520_ _04529_ _04530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_36_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08441_ _03918_ _00415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05653_ soc.cpu.ALU.ny _01561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_1_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_210_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_184_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_229_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08372_ soc.spi_video_ram_1.write_fifo.fifo_mem\[26\]\[14\] _02246_ _03877_ _03882_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_189_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05584_ _01490_ _01491_ _01492_ _01493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_07323_ _02926_ soc.spi_video_ram_1.write_fifo.fifo_mem\[15\]\[28\] _02722_ _02973_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_123_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07254_ soc.spi_video_ram_1.write_fifo.fifo_mem\[16\]\[9\] soc.spi_video_ram_1.write_fifo.fifo_mem\[17\]\[9\]
+ soc.spi_video_ram_1.write_fifo.fifo_mem\[18\]\[9\] soc.spi_video_ram_1.write_fifo.fifo_mem\[19\]\[9\]
+ _02903_ _02904_ _02905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_191_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06205_ soc.spi_video_ram_1.buffer_index\[4\] _02090_ _02091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_07185_ soc.spi_video_ram_1.write_fifo.fifo_mem\[12\]\[6\] soc.spi_video_ram_1.write_fifo.fifo_mem\[13\]\[6\]
+ soc.spi_video_ram_1.write_fifo.fifo_mem\[14\]\[6\] soc.spi_video_ram_1.write_fifo.fifo_mem\[15\]\[6\]
+ _02680_ _02838_ _02839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_121_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_219_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_180_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06136_ _02028_ _01962_ _02029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_2_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06067_ _01950_ _01959_ _01960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_236_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09826_ _04741_ _04753_ _04754_ _04755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_24_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09757_ _04695_ _04708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
Xclkbuf_leaf_5_wb_clk_i clknet_5_0_0_wb_clk_i clknet_leaf_5_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_06969_ _01428_ soc.spi_video_ram_1.current_state\[0\] _02630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_210_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2104 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08708_ _03511_ _04046_ _04064_ _00536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_2115 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2126 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09688_ soc.cpu.PC.REG.data\[8\] soc.rom_loader.current_address\[8\] _04638_ _04660_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_2137 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_271_wb_clk_i clknet_5_6_0_wb_clk_i clknet_leaf_271_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_2148 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2159 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08639_ _04024_ _00507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_242_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_200_wb_clk_i clknet_5_19_0_wb_clk_i clknet_leaf_200_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_214_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11650_ _00711_ clknet_leaf_28_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[20\]\[18\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_230_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_35_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10601_ _05277_ _05278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_208_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11581_ _00647_ clknet_leaf_26_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[22\]\[17\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xfanout85 soc.cpu.AReg.clk net85 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_10532_ soc.ram_encoder_0.address\[7\] soc.cpu.AReg.data\[7\] _05227_ _05236_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_122_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_221_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_13_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_167_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10463_ _05171_ _05184_ _05185_ _01170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_109_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_202_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_164_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_104_1594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12202_ _01230_ clknet_leaf_40_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[19\]\[13\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_136_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10394_ _02244_ soc.spi_video_ram_1.write_fifo.fifo_mem\[6\]\[13\] _05135_ _05139_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_89_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_139_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12133_ _01161_ clknet_leaf_289_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[6\]\[25\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_85_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12064_ _01107_ clknet_leaf_112_wb_clk_i soc.rom_loader.current_address\[4\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_46_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11015_ _00081_ clknet_leaf_42_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[16\]\[11\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_93_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_238_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4040 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_213_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4051 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_237_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4062 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_218_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4073 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4084 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4095 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_234_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11917_ _00976_ clknet_leaf_122_wb_clk_i soc.cpu.instruction\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_185_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_233_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2693 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11848_ _00907_ clknet_leaf_122_wb_clk_i soc.rom_encoder_0.request_data_out\[9\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_21_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1970 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_226_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1981 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1992 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_1314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11779_ _00840_ clknet_leaf_104_wb_clk_i soc.rom_encoder_0.output_buffer\[10\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_109_1483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_220_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_147_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_75_wb_clk_i clknet_5_8_0_wb_clk_i clknet_leaf_75_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_103_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08990_ _04217_ _00665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_86_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07941_ soc.spi_video_ram_1.write_fifo.fifo_mem\[4\]\[20\] soc.spi_video_ram_1.write_fifo.fifo_mem\[5\]\[20\]
+ soc.spi_video_ram_1.write_fifo.fifo_mem\[6\]\[20\] soc.spi_video_ram_1.write_fifo.fifo_mem\[7\]\[20\]
+ _02764_ _02723_ _03583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_102_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_190_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07872_ _02704_ soc.spi_video_ram_1.write_fifo.fifo_mem\[11\]\[22\] _02578_ _03516_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_99_1405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09611_ soc.rom_encoder_0.input_buffer\[11\] _04609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_28_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_214_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06823_ _02484_ _02481_ _02499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_83_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_237_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06754_ soc.rom_encoder_0.current_state\[0\] _02433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
X_09542_ _01403_ _04558_ _04561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_110_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05705_ _01585_ _01597_ _01608_ _01611_ _01612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_77_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06685_ _02392_ _00186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09473_ _01437_ _01417_ _02624_ _04517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_224_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08424_ _03909_ _00407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_93_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05636_ soc.spi_video_ram_1.output_buffer\[2\] soc.spi_video_ram_1.output_buffer\[3\]
+ _01467_ _01545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_244_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_145_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_205_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_212_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08355_ soc.spi_video_ram_1.write_fifo.fifo_mem\[26\]\[6\] _02403_ _03866_ _03873_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_127_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05567_ soc.spi_video_ram_1.buffer_index\[1\] _01475_ _01476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_205_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07306_ _02612_ soc.spi_video_ram_1.write_fifo.fifo_mem\[21\]\[10\] _02956_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__and2_1
X_08286_ _03835_ _00343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_149_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05498_ soc.spi_video_ram_1.initialized soc.spi_video_ram_1.current_state\[2\] _01413_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07237_ soc.spi_video_ram_1.write_fifo.fifo_mem\[0\]\[9\] soc.spi_video_ram_1.write_fifo.fifo_mem\[1\]\[9\]
+ soc.spi_video_ram_1.write_fifo.fifo_mem\[2\]\[9\] soc.spi_video_ram_1.write_fifo.fifo_mem\[3\]\[9\]
+ _02680_ _02722_ _02888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_165_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_203_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_146_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_192_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07168_ _02822_ _00238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_106_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06119_ _01969_ _02012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_1_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07099_ _02678_ _02749_ _02755_ _02586_ _02756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_156_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_232_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09809_ _04739_ _04740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_8_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_219_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_216_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_243_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11702_ _00763_ clknet_leaf_200_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[9\]\[4\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_215_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_231_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11633_ _00694_ clknet_leaf_216_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[20\]\[1\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_243_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_202_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_196_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_180_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11564_ _00630_ clknet_leaf_205_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[22\]\[0\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_106_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10515_ _05221_ _05224_ _05226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11495_ _00561_ clknet_leaf_23_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[24\]\[18\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_137_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10446_ _02053_ _05173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xcaravel_hack_soc_130 la_data_out[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xcaravel_hack_soc_141 la_data_out[13] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_137_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xcaravel_hack_soc_152 la_data_out[24] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_108_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xcaravel_hack_soc_163 la_data_out[36] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_48_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xcaravel_hack_soc_174 la_data_out[47] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xcaravel_hack_soc_185 la_data_out[58] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_10377_ _02227_ soc.spi_video_ram_1.write_fifo.fifo_mem\[6\]\[5\] _05124_ _05130_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xcaravel_hack_soc_196 wbs_dat_o[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_124_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12116_ _01144_ clknet_leaf_244_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[6\]\[8\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12047_ net24 clknet_leaf_95_wb_clk_i soc.rom_encoder_0.data_out\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_46_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_211_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_193_wb_clk_i clknet_5_28_0_wb_clk_i clknet_leaf_193_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_187_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_37_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_219_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_122_wb_clk_i clknet_5_15_0_wb_clk_i clknet_leaf_122_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_20_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_241_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3180 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_206_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_209_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_1357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06470_ soc.spi_video_ram_1.write_fifo.fifo_mem\[16\]\[25\] _02268_ _02216_ _02269_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_59_1488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_107_1409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_221_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08140_ _03735_ _00297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_109_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_222_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_186_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08071_ soc.spi_video_ram_1.write_fifo.fifo_mem\[11\]\[13\] _02244_ _03691_ _03695_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_147_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07022_ _02680_ _02681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_174_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_196_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08973_ soc.spi_video_ram_1.write_fifo.fifo_mem\[22\]\[28\] _02353_ _04177_ _04208_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_25_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07924_ _02931_ _03566_ _03567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_4809 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_233_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_131_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_29_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07855_ _03481_ _03489_ _03498_ _02567_ _03499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_112_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_29_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06806_ soc.ram_encoder_0.current_state\[0\] _02482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_07786_ soc.spi_video_ram_1.write_fifo.fifo_mem\[23\]\[23\] _03431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_84_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_227_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09525_ _01836_ _01993_ _02058_ _04548_ _04549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_65_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_231_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06737_ _02424_ _00206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_225_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_164_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xclkbuf_3_5_0_wb_clk_i clknet_2_2_0_wb_clk_i clknet_3_5_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_196_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09456_ _03770_ _04473_ _04503_ _00846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XPHY_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_06668_ _02167_ soc.spi_video_ram_1.write_fifo.fifo_mem\[12\]\[23\] _02356_ _02382_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_80_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_213_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_101_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05619_ soc.spi_video_ram_1.output_buffer\[22\] soc.spi_video_ram_1.output_buffer\[23\]
+ _01468_ _01528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_08407_ soc.spi_video_ram_1.write_fifo.fifo_mem\[27\]\[1\] _02393_ _03899_ _03901_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_51_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_71_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06599_ _02344_ _00148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09387_ net69 _04430_ _04433_ _04451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_184_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08338_ soc.spi_video_ram_1.write_fifo.write_pointer\[2\] _03862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_240_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_162_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_201_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08269_ _02558_ _03823_ _03824_ _00337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_10300_ soc.rom_loader.current_address\[6\] _05082_ _05084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_153_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_193_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11280_ _00346_ clknet_leaf_213_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[1\]\[6\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_119_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_175_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10231_ _02240_ soc.spi_video_ram_1.write_fifo.fifo_mem\[5\]\[11\] _05041_ _05043_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_156_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_238_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10162_ _01381_ _04997_ _01057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_156_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10093_ _04928_ _04943_ _04944_ _04945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_134_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_16_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_75_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_223_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10995_ _00061_ clknet_leaf_264_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[17\]\[20\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_188_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_206_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_167_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_203_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11616_ _00682_ clknet_leaf_241_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[21\]\[23\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_180_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_223_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11547_ _00613_ clknet_leaf_319_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[25\]\[12\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_184_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11478_ _00544_ clknet_leaf_180_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[24\]\[1\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10429_ net90 _05017_ _05156_ _01165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_125_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_217_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_125_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_154_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_170_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_303_wb_clk_i clknet_5_4_0_wb_clk_i clknet_leaf_303_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05970_ soc.video_generator_1.v_count\[8\] soc.video_generator_1.v_count\[7\] _01849_
+ soc.video_generator_1.v_count\[5\] _01863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_140_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_152_1451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_238_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07640_ _02695_ soc.spi_video_ram_1.write_fifo.fifo_mem\[16\]\[14\] _03286_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_20_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07571_ _03021_ soc.spi_video_ram_1.write_fifo.fifo_mem\[13\]\[13\] _03217_ _03024_
+ _03218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_213_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_207_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09310_ _04405_ _00797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06522_ _02157_ soc.spi_video_ram_1.write_fifo.fifo_mem\[0\]\[18\] _02290_ _02299_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_178_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_228_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09241_ _04368_ _00765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06453_ _02257_ _00089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_194_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_146_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09172_ _04317_ _04326_ _04327_ _00737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_06384_ _02210_ _00067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_119_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_193_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08123_ soc.video_generator_1.h_count\[7\] _03723_ _03724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_190_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08054_ soc.spi_video_ram_1.write_fifo.fifo_mem\[11\]\[5\] _02401_ _03680_ _03686_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_07005_ _02650_ _02664_ _02618_ _02665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_116_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_227_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_227_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_157_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_6008 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_89_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6019 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08956_ _04199_ _00649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_4606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07907_ _02920_ soc.spi_video_ram_1.write_fifo.fifo_mem\[17\]\[21\] _03550_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_4639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3905 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_56_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08887_ _04162_ _00617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_84_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3916 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3927 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3938 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07838_ soc.spi_video_ram_1.write_fifo.fifo_mem\[23\]\[22\] _03482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_3949 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_205_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07769_ _02831_ _03407_ _03413_ _03414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_25_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09508_ _02262_ soc.cpu.AReg.data\[6\] _04339_ _04539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XPHY_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_197_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10780_ _03246_ _05358_ _05373_ _01300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_40_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_207_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_158_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_73_1249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09439_ soc.rom_encoder_0.request_data_out\[5\] _03767_ _04490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XPHY_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_129_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_185_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11401_ _00467_ clknet_leaf_14_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[2\]\[11\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_122_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_166_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_197_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11332_ _00398_ clknet_leaf_186_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[27\]\[0\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_125_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_177_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_180_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_158_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11263_ _00329_ clknet_leaf_151_wb_clk_i soc.ram_encoder_0.output_buffer\[9\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_137_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_218_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10214_ _02223_ soc.spi_video_ram_1.write_fifo.fifo_mem\[5\]\[3\] _05030_ _05034_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_11194_ _00260_ clknet_leaf_196_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[11\]\[4\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_6520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_171_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_171_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10145_ soc.ram_data_out\[15\] _04928_ _04984_ _04985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_79_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_6564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5830 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_212_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5841 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5852 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5863 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10076_ soc.ram_encoder_0.request_data_out\[0\] _04930_ _04931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_5874 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_5885 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5896 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_130_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_236_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_225_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_95_1474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10978_ _00044_ clknet_leaf_140_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[17\]\[3\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_147_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_169_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_172_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08810_ _04121_ _00581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_113_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09790_ _02270_ soc.spi_video_ram_1.write_fifo.fifo_mem\[3\]\[26\] _04696_ _04725_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_234_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08741_ soc.spi_video_ram_1.write_fifo.fifo_mem\[24\]\[7\] _02405_ _04076_ _04084_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_05953_ _01842_ _01845_ _01846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_152_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05884_ _01595_ _01779_ _01780_ soc.cpu.PC.in\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_08672_ soc.spi_video_ram_1.write_fifo.fifo_mem\[15\]\[9\] _02409_ _04032_ _04042_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_66_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_187_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_242_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07623_ soc.spi_video_ram_1.write_fifo.fifo_mem\[15\]\[25\] _03270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_54_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_35_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07554_ _02924_ soc.spi_video_ram_1.write_fifo.fifo_mem\[30\]\[13\] _03200_ _02908_
+ _03201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_74_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06505_ _02277_ _02290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_07485_ _02645_ soc.spi_video_ram_1.write_fifo.fifo_mem\[6\]\[12\] _03132_ _02577_
+ _03133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_195_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_167_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09224_ _02179_ _03729_ _04358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06436_ soc.spi_video_ram_1.fifo_in_data\[14\] _02246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_33_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_202_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09155_ _01931_ soc.video_generator_1.v_count\[1\] _01866_ _04315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_06367_ _02157_ soc.spi_video_ram_1.write_fifo.fifo_mem\[17\]\[18\] _02193_ _02202_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_163_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_1413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08106_ soc.display_clks_before_active\[0\] _03713_ _00285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_175_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_296_wb_clk_i clknet_5_4_0_wb_clk_i clknet_leaf_296_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_107_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_194_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_162_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09086_ _04273_ _00705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06298_ _02160_ _00031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_102_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08037_ _03665_ _03674_ _03675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_135_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_5_26_0_wb_clk_i clknet_4_13_0_wb_clk_i clknet_5_26_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_27_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5104 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_231_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5115 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5126 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09988_ _04833_ _04876_ _04877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_5137 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_213_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5148 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_190_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5159 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_236_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08939_ soc.spi_video_ram_1.write_fifo.fifo_mem\[22\]\[11\] _02414_ _04189_ _04191_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_4425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_170_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3702 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3713 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11950_ _01009_ clknet_leaf_156_wb_clk_i soc.ram_encoder_0.request_data_out\[3\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3724 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3735 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3746 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_218_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3757 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10901_ soc.spi_video_ram_1.write_fifo.fifo_mem\[8\]\[7\] soc.spi_video_ram_1.fifo_in_data\[7\]
+ _05431_ _05439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_3768 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_229_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3779 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11881_ _00940_ clknet_5_19_0_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[3\]\[7\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_232_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10832_ _02258_ soc.spi_video_ram_1.write_fifo.fifo_mem\[7\]\[20\] _05389_ _05402_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_246_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_201_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_158_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10763_ soc.spi_video_ram_1.write_fifo.fifo_mem\[31\]\[17\] soc.spi_video_ram_1.fifo_in_address\[1\]
+ _05355_ _05365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_13_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_157_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10694_ soc.spi_video_ram_1.fifo_in_data\[14\] _05325_ _05328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_12_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_154_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_240_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11315_ _00381_ clknet_leaf_1_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[26\]\[12\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_114_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12295_ _01323_ clknet_leaf_73_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[7\]\[19\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_218_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11246_ _00312_ clknet_leaf_24_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[10\]\[17\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_64_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_190_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11177_ _00243_ clknet_leaf_60_wb_clk_i soc.spi_video_ram_1.output_buffer\[13\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_6361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_132_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_7_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10128_ _04863_ _04947_ _04948_ _04971_ _04972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_6394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_231_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_5682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5693 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10059_ soc.ram_encoder_0.initializing_step\[4\] soc.ram_encoder_0.initializing_step\[2\]
+ _04916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_76_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4970 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_235_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_224_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4981 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_29_wb_clk_i clknet_5_9_0_wb_clk_i clknet_leaf_29_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_4992 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07270_ _02919_ _02920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_177_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_176_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06221_ _02087_ _02101_ _02106_ _02094_ _02107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_192_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06152_ _01972_ _01973_ _02044_ _01925_ _02045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_144_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06083_ _01907_ _01975_ _01976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_160_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09911_ _04818_ _04819_ _04553_ _04820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_67_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_217_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09842_ soc.cpu.instruction\[5\] _04740_ _04767_ _04768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_59_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_140_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_218_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09773_ _04716_ _00950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06985_ _02644_ _02645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XTAP_3009 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_132_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08724_ soc.spi_video_ram_1.write_fifo.write_pointer\[1\] _01405_ _03863_ _04074_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_113_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05936_ _01826_ _01830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_41_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08655_ _04033_ _00514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_214_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05867_ _01586_ _01758_ _01761_ _01765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_42_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07606_ _02901_ _03245_ _03252_ _02970_ _03253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_1618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08586_ _02175_ soc.spi_video_ram_1.write_fifo.fifo_mem\[2\]\[27\] _03966_ _03996_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_241_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_230_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05798_ _01553_ _01615_ soc.cpu.AReg.data\[6\] _01592_ _01700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_35_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07537_ _03146_ _03184_ _03185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_224_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_210_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07468_ _02901_ _03108_ _03115_ _02910_ _03116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_168_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_139_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_194_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09207_ _00011_ _01713_ _04349_ _00750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06419_ _02234_ _00078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07399_ _03047_ soc.spi_video_ram_1.write_fifo.fifo_mem\[10\]\[11\] _03048_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_176_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09138_ _04294_ _04302_ _04303_ _00727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_163_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_151_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09069_ _04264_ _00697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_190_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11100_ _00166_ clknet_leaf_202_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[12\]\[9\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12080_ soc.cpu.PC.in\[3\] net84 soc.cpu.AReg.data\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_235_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11031_ _00097_ clknet_leaf_271_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[16\]\[27\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_85_1495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_215_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_172_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_237_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_44_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_4233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_217_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_206_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11933_ _00992_ clknet_leaf_165_wb_clk_i soc.ram_encoder_0.input_bits_left\[4\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_73_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2820 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_233_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2831 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2842 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2853 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11864_ _00923_ clknet_leaf_109_wb_clk_i soc.rom_encoder_0.request_address\[9\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_17_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2864 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2875 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_127_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2886 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_242_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_183_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10815_ _05377_ _05393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_2897 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11795_ _00011_ clknet_leaf_132_wb_clk_i soc.spi_video_ram_1.fifo_write_request vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_246_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_207_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10746_ _05343_ _05355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_159_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_147_wb_clk_i clknet_5_28_0_wb_clk_i clknet_leaf_147_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_70_1753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10677_ _02231_ soc.spi_video_ram_1.write_fifo.fifo_mem\[29\]\[7\] _05310_ _05318_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_199_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_177_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12347_ _01375_ clknet_leaf_287_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[8\]\[26\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_154_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_142_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_5_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12278_ _01306_ clknet_leaf_265_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[7\]\[2\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_190_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11229_ _00295_ clknet_leaf_191_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[10\]\[0\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_136_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_229_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_214_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6180 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_136_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06770_ soc.rom_encoder_0.initializing_step\[4\] soc.rom_encoder_0.initializing_step\[3\]
+ soc.rom_encoder_0.initializing_step\[2\] soc.rom_encoder_0.initializing_step\[1\]
+ _02449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_82_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_95_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_188_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05721_ _01617_ _01626_ _01627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_64_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08440_ soc.spi_video_ram_1.write_fifo.fifo_mem\[27\]\[17\] _02337_ _03910_ _03918_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_05652_ _01557_ _01559_ _01560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_24_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_223_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_212_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08371_ _03881_ _00382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05583_ _01462_ _01485_ _01492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_225_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07322_ _02971_ soc.spi_video_ram_1.write_fifo.fifo_mem\[14\]\[28\] _02972_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_143_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_182_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_176_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07253_ _02894_ _02904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_104_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_192_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06204_ _01464_ _01494_ _02090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07184_ _02646_ _02838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_69_1413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06135_ _01945_ _01958_ _01960_ _02028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_117_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_238_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_191_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_160_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06066_ soc.video_generator_1.h_count\[8\] _01838_ soc.video_generator_1.h_count\[9\]
+ _01959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
XFILLER_28_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_232_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_235_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_160_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09825_ net7 _04566_ _04754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_150_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_219_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_246_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09756_ _04707_ _00942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06968_ _02624_ _02629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_27_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08707_ _04063_ _04048_ _04064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05919_ _01811_ _01814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_2105 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09687_ _04618_ _04658_ _04659_ _00921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_2116 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06899_ soc.ram_encoder_0.request_address\[1\] _02506_ _02562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_64_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2127 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_215_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2138 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2149 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08638_ _02165_ soc.spi_video_ram_1.write_fifo.fifo_mem\[30\]\[22\] _03999_ _04024_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_82_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_199_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_243_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08569_ _03987_ _00474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_180_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10600_ _05276_ _05277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_211_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11580_ _00646_ clknet_leaf_26_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[22\]\[16\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_161_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout86 soc.cpu.AReg.clk net86 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_195_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10531_ _05235_ _01189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xclkbuf_leaf_240_wb_clk_i clknet_5_17_0_wb_clk_i clknet_leaf_240_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_11_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_122_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10462_ soc.cpu.PC.in\[4\] _05172_ _05173_ _05185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_108_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12201_ _01229_ clknet_leaf_2_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[19\]\[12\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_202_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_178_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10393_ _05138_ _01148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_191_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12132_ _01160_ clknet_leaf_301_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[6\]\[24\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_97_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_12063_ _01106_ clknet_leaf_112_wb_clk_i soc.rom_loader.current_address\[3\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_2_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_145_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_215_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11014_ _00080_ clknet_leaf_13_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[16\]\[10\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_78_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4030 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4041 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4052 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_77_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4063 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4074 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4085 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4096 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11916_ _00975_ clknet_leaf_119_wb_clk_i soc.cpu.instruction\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_46_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_205_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11847_ _00906_ clknet_leaf_169_wb_clk_i soc.rom_encoder_0.request_data_out\[8\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2694 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1960 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1971 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1982 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1993 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11778_ _00839_ clknet_leaf_93_wb_clk_i soc.rom_encoder_0.output_buffer\[9\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_109_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_222_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_147_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_201_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_1495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10729_ _05346_ _01276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_105_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_220_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_196_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_157_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_154_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_4_7_0_wb_clk_i clknet_3_3_0_wb_clk_i clknet_4_7_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_157_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07940_ _02768_ _03581_ _03582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_218_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_233_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_44_wb_clk_i clknet_5_6_0_wb_clk_i clknet_leaf_44_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_155_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07871_ _02689_ soc.spi_video_ram_1.write_fifo.fifo_mem\[10\]\[22\] _03515_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09610_ _04607_ _04586_ _04608_ _00895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_228_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06822_ _02491_ _02485_ _02498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_42_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09541_ _01446_ _04552_ _02312_ _04560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06753_ _02432_ _00214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_83_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05704_ _01585_ _01610_ _01611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_52_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09472_ _02542_ _04515_ _04516_ _00849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_24_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06684_ soc.spi_video_ram_1.write_fifo.fifo_mem\[14\]\[0\] _02310_ _02391_ _02392_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_36_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_184_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08423_ soc.spi_video_ram_1.write_fifo.fifo_mem\[27\]\[9\] _02409_ _03899_ _03909_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_24_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05635_ _01470_ _01543_ _01544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_240_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_1483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08354_ _03872_ _00374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05566_ _01460_ _01474_ _01464_ _01475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_138_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07305_ _02696_ soc.spi_video_ram_1.write_fifo.fifo_mem\[23\]\[10\] _02895_ _02955_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08285_ _02126_ soc.spi_video_ram_1.write_fifo.fifo_mem\[1\]\[3\] _03831_ _03835_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_05497_ soc.spi_video_ram_1.current_state\[0\] _01408_ _01411_ _01412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_07236_ _02589_ _02886_ _02640_ _02887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_118_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07167_ soc.spi_video_ram_1.output_buffer\[18\] _02821_ _02633_ _02822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_106_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06118_ _01922_ _02009_ _02010_ _02011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_246_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_79_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07098_ _02750_ _02751_ _02754_ _02693_ _02643_ _02755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_105_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_160_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06049_ _01932_ _01941_ _01942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_132_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_1487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09808_ _02434_ _02435_ _04738_ _04739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_60_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_210_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09739_ _02219_ soc.spi_video_ram_1.write_fifo.fifo_mem\[3\]\[1\] _04697_ _04699_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_21_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_242_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11701_ _00762_ clknet_leaf_198_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[9\]\[3\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_152_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_230_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11632_ _00693_ clknet_leaf_207_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[20\]\[0\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_208_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11563_ _00629_ clknet_leaf_297_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[25\]\[28\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_156_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_156_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_221_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10514_ _05222_ _05225_ _01182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_109_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11494_ _00560_ clknet_leaf_19_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[24\]\[17\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_109_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xcaravel_hack_soc_120 io_out[26] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_10445_ _05170_ _05172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_155_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xcaravel_hack_soc_131 la_data_out[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_100_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xcaravel_hack_soc_142 la_data_out[14] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_139_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xcaravel_hack_soc_153 la_data_out[25] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xcaravel_hack_soc_164 la_data_out[37] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xcaravel_hack_soc_175 la_data_out[48] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xcaravel_hack_soc_186 la_data_out[59] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_3_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10376_ _05129_ _01140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_237_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xcaravel_hack_soc_197 wbs_dat_o[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_12115_ _01143_ clknet_leaf_243_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[6\]\[7\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_69_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_219_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_151_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12046_ net23 clknet_5_31_0_wb_clk_i soc.rom_encoder_0.data_out\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_133_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_238_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_4_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_234_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_opt_2_0_wb_clk_i clknet_5_11_0_wb_clk_i clknet_opt_2_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_34_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3170 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3181 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_162_wb_clk_i clknet_5_27_0_wb_clk_i clknet_leaf_162_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_185_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_233_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_222_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_226_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1790 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_187_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08070_ _03694_ _00268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07021_ _02679_ _02680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_200_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_192_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_118_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08972_ _04207_ _00657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_115_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07923_ soc.spi_video_ram_1.write_fifo.fifo_mem\[31\]\[21\] _03566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_190_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_29_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07854_ _02767_ _03490_ _03497_ _02970_ _03498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_57_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_229_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06805_ soc.ram_encoder_0.current_state\[1\] _02481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_84_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07785_ _02693_ _03426_ _03429_ _02901_ _03430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_09524_ soc.video_generator_1.h_count\[6\] _04546_ _04547_ _04548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_71_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06736_ soc.spi_video_ram_1.write_fifo.fifo_mem\[14\]\[20\] _02343_ _02390_ _02424_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_37_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_224_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09455_ _02461_ _02541_ _04502_ _04503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XPHY_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_06667_ _02381_ _00179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_51_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08406_ _03900_ _00398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_212_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05618_ _01463_ _01526_ _01527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_75_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09386_ net69 _04430_ _04448_ _00828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_06598_ soc.spi_video_ram_1.write_fifo.fifo_mem\[13\]\[20\] _02343_ _02316_ _02344_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_123_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_196_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08337_ _03861_ _00368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_178_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05549_ _01458_ _01459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_229_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08268_ soc.ram_encoder_0.output_buffer\[17\] _02555_ _03824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_20_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_203_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07219_ soc.spi_video_ram_1.write_fifo.fifo_mem\[28\]\[8\] soc.spi_video_ram_1.write_fifo.fifo_mem\[29\]\[8\]
+ soc.spi_video_ram_1.write_fifo.fifo_mem\[30\]\[8\] soc.spi_video_ram_1.write_fifo.fifo_mem\[31\]\[8\]
+ _02607_ _02636_ _02871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_158_1319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_192_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08199_ soc.rom_encoder_0.output_buffer\[16\] _03766_ _03767_ soc.rom_encoder_0.request_data_out\[12\]
+ _03768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_88_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10230_ _05042_ _01081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_69_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10161_ _02481_ _04993_ _04994_ _02510_ _04997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_161_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_216_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10092_ net4 _04834_ _04944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_48_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_216_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10994_ _00060_ clknet_leaf_68_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[17\]\[19\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_243_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_1509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_215_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_204_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_16_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_71_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_231_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_70_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_243_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11615_ _00681_ clknet_leaf_250_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[21\]\[22\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_54_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11546_ _00612_ clknet_leaf_33_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[25\]\[11\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_11_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_204_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11477_ _00543_ clknet_leaf_187_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[24\]\[0\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_137_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10428_ net90 _01181_ _05156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_178_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10359_ _01819_ _05104_ _05119_ _01133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_234_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_183_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_191_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_239_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_12029_ _01088_ clknet_leaf_67_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[5\]\[17\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_78_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07570_ _02919_ soc.spi_video_ram_1.write_fifo.fifo_mem\[12\]\[13\] _03217_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_53_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_206_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06521_ _02298_ _00116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_185_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09240_ _02229_ soc.spi_video_ram_1.write_fifo.fifo_mem\[9\]\[6\] _04365_ _04368_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06452_ soc.spi_video_ram_1.write_fifo.fifo_mem\[16\]\[19\] _02256_ _02238_ _02257_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_72_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_221_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_178_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09171_ _02034_ _04325_ _04327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_33_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06383_ _02173_ soc.spi_video_ram_1.write_fifo.fifo_mem\[17\]\[26\] _02181_ _02210_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_08122_ _03713_ _03722_ _03723_ _00291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_222_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_190_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08053_ _03685_ _00260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_119_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07004_ soc.spi_video_ram_1.write_fifo.fifo_mem\[20\]\[1\] soc.spi_video_ram_1.write_fifo.fifo_mem\[21\]\[1\]
+ soc.spi_video_ram_1.write_fifo.fifo_mem\[22\]\[1\] soc.spi_video_ram_1.write_fifo.fifo_mem\[23\]\[1\]
+ _02651_ _02593_ _02664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_157_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_190_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6009 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_5_16_0_wb_clk_i clknet_4_8_0_wb_clk_i clknet_5_16_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_116_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08955_ soc.spi_video_ram_1.write_fifo.fifo_mem\[22\]\[19\] _02341_ _04189_ _04199_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_4607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_233_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07906_ soc.spi_video_ram_1.write_fifo.fifo_mem\[18\]\[21\] soc.spi_video_ram_1.write_fifo.fifo_mem\[19\]\[21\]
+ _02651_ _03549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_57_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_243_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08886_ soc.spi_video_ram_1.write_fifo.fifo_mem\[25\]\[16\] _02335_ _04155_ _04162_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_170_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3906 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3917 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3928 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07837_ _02693_ _03477_ _03480_ _02707_ _03481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XTAP_3939 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_99_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_246_1612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07768_ _03408_ _03409_ _03412_ _02976_ _02929_ _03413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_244_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_225_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09507_ _04538_ _00862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_164_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06719_ _02415_ _00197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_73_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07699_ _02573_ _03344_ _03345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_72_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_1682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_188_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09438_ _04473_ _04488_ _04489_ _00842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_213_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_184_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_199_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09369_ _04439_ _04440_ _00821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_197_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_240_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_201_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11400_ _00466_ clknet_leaf_18_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[2\]\[10\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_162_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_166_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_138_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11331_ _00397_ clknet_leaf_298_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[26\]\[28\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_10_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_123_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11262_ _00328_ clknet_leaf_151_wb_clk_i soc.ram_encoder_0.output_buffer\[8\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_49_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_238_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10213_ _05033_ _01073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_106_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_6510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11193_ _00259_ clknet_leaf_260_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[11\]\[3\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_6521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10144_ _04871_ _04930_ _04926_ _04983_ _04984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_6554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5820 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5831 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5842 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_88_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5853 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_114_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10075_ _04929_ _04930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_153_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5864 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5875 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5886 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5897 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_212_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_186_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10977_ _00043_ clknet_leaf_197_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[17\]\[2\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_108_1505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_203_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_176_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_50_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_12_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_223_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_200_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_190_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11529_ _00595_ clknet_leaf_243_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[23\]\[23\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_156_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_217_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_61_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08740_ _04083_ _00549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_113_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05952_ soc.video_generator_1.h_count\[5\] soc.video_generator_1.h_count\[6\] _01845_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_230_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_238_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08671_ _04041_ _00522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05883_ _01552_ soc.cpu.ALU.zx soc.cpu.AReg.data\[11\] _01591_ _01780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_66_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07622_ _03264_ _03265_ _03268_ _02691_ _02929_ _03269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_96_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_199_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_226_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_207_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07553_ _02907_ _03199_ _03200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_165_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_146_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06504_ _02289_ _00108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_228_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07484_ _02919_ _03131_ _03132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_146_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09223_ _04341_ _02539_ _04357_ _00758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_166_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06435_ _02245_ _00083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_179_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_241_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09154_ _01860_ soc.video_generator_1.v_count\[8\] soc.video_generator_1.v_count\[7\]
+ _01849_ _04314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
X_06366_ _02201_ _00058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_33_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_163_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08105_ _01959_ _03712_ _01380_ _03713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_4
X_09085_ _02145_ soc.spi_video_ram_1.write_fifo.fifo_mem\[20\]\[12\] _04270_ _04273_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06297_ _02159_ soc.spi_video_ram_1.write_fifo.fifo_mem\[18\]\[19\] _02141_ _02160_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_163_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08036_ _03667_ _03669_ _03671_ _03673_ _02568_ _03674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_163_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_239_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5105 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_265_wb_clk_i clknet_5_7_0_wb_clk_i clknet_leaf_265_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_192_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5116 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09987_ _04874_ _04875_ _04876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_27_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_5127 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5138 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5149 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08938_ _04190_ _00640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_4415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3703 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08869_ soc.spi_video_ram_1.write_fifo.fifo_mem\[25\]\[8\] _02407_ _04144_ _04153_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_3714 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_213_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3725 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3736 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3747 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10900_ _05438_ _01355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3758 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11880_ _00939_ clknet_leaf_247_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[3\]\[6\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3769 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_189_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10831_ _05401_ _01323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_246_1442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_26_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_73_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_207_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_183_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10762_ _05364_ _01291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_25_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_232_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_186_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_160_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_240_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_185_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10693_ _03202_ _05324_ _05327_ _01259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_139_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_154_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_4_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11314_ _00380_ clknet_leaf_34_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[26\]\[11\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12294_ _01322_ clknet_leaf_80_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[7\]\[18\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_154_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11245_ _00311_ clknet_leaf_25_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[10\]\[16\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_107_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_175_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_79_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11176_ _00242_ clknet_leaf_56_wb_clk_i soc.spi_video_ram_1.output_buffer\[14\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_6351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_218_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_171_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10127_ soc.ram_encoder_0.request_data_out\[11\] _04929_ _04971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_6384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10058_ soc.ram_encoder_0.initialized _04254_ _04915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_57_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5694 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_7_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4960 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_4971 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4982 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_236_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4993 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_208_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_69_wb_clk_i clknet_5_11_0_wb_clk_i clknet_leaf_69_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_189_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_232_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06220_ _02091_ _02102_ _02105_ _02087_ _02106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_176_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_191_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06151_ _01977_ _02043_ _02044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_8_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06082_ _01893_ _01894_ _01899_ _01975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_171_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09910_ soc.rom_encoder_0.initializing_step\[1\] _02459_ _03763_ _02460_ _04819_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_160_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09841_ _04588_ _04761_ _04762_ _04766_ _04767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_98_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09772_ _02252_ soc.spi_video_ram_1.write_fifo.fifo_mem\[3\]\[17\] _04708_ _04716_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06984_ _02572_ _02644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XTAP_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08723_ _04073_ _00542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_67_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05935_ _01805_ _01798_ _01811_ _01829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_239_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_187_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08654_ soc.spi_video_ram_1.write_fifo.fifo_mem\[15\]\[0\] _02310_ _04032_ _04033_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_242_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05866_ _01762_ _01754_ _01756_ _01764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_54_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_96_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07605_ _02588_ _03248_ _03251_ _03252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_1608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_208_1702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08585_ _03995_ _00482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05797_ _01615_ _01698_ _01699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_74_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07536_ _02620_ _03165_ _03183_ _03019_ _03184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_74_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_208_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_222_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_167_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07467_ _02642_ _03111_ _03114_ _03115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_126_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_161_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09206_ soc.spi_video_ram_1.fifo_in_data\[7\] _04346_ _04349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_202_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06418_ soc.spi_video_ram_1.write_fifo.fifo_mem\[16\]\[8\] _02233_ _02217_ _02234_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_33_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_10_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07398_ _02783_ _03047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_210_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09137_ soc.spi_video_ram_1.state_counter\[5\] _04300_ _04303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06349_ _02192_ _00050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_87_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_108_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_194_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_163_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09068_ _02225_ soc.spi_video_ram_1.write_fifo.fifo_mem\[20\]\[4\] _04259_ _04264_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_237_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_150_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08019_ soc.spi_video_ram_1.write_fifo.fifo_mem\[0\]\[16\] soc.spi_video_ram_1.write_fifo.fifo_mem\[1\]\[16\]
+ soc.spi_video_ram_1.write_fifo.fifo_mem\[2\]\[16\] soc.spi_video_ram_1.write_fifo.fifo_mem\[3\]\[16\]
+ _02701_ _02737_ _03657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_215_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_11030_ _00096_ clknet_leaf_287_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[16\]\[26\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_46_1447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_137_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_4245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_218_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11932_ _00991_ clknet_leaf_164_wb_clk_i soc.ram_encoder_0.input_bits_left\[3\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_4289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2810 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2821 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_232_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2832 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_5_9_0_wb_clk_i clknet_4_4_0_wb_clk_i clknet_5_9_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XTAP_3577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2843 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11863_ _00922_ clknet_leaf_105_wb_clk_i soc.rom_encoder_0.request_address\[8\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_79_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2854 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2865 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2876 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10814_ _05389_ _05392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_2887 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2898 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_220_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_214_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11794_ _00855_ clknet_5_24_0_wb_clk_i soc.spi_video_ram_1.buffer_index\[5\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_246_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10745_ _05354_ _01284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_40_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_146_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10676_ _05317_ _01252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_224_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_167_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_12346_ _01374_ clknet_leaf_237_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[8\]\[25\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_154_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_153_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_187_wb_clk_i clknet_5_29_0_wb_clk_i clknet_leaf_187_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_245_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_142_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12277_ _01305_ clknet_leaf_245_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[7\]\[1\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_9_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_64_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11228_ _00294_ clknet_leaf_86_wb_clk_i soc.video_generator_1.h_count\[9\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_2
XTAP_6170 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11159_ _00225_ clknet_leaf_105_wb_clk_i soc.rom_encoder_0.output_buffer\[4\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_96_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_190_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6181 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_191_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_49_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_5480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05720_ _01561_ _01625_ _01626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_23_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_224_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_237_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4790 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_184_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05651_ _01558_ soc.cpu.ALU.x\[0\] _01559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_75_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08370_ soc.spi_video_ram_1.write_fifo.fifo_mem\[26\]\[13\] _02244_ _03877_ _03881_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_56_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05582_ soc.spi_video_ram_1.output_buffer\[9\] soc.spi_video_ram_1.output_buffer\[8\]
+ _01461_ _01491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_177_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07321_ _02574_ _02971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_108_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_177_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_204_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_149_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_221_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_242_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07252_ _02902_ _02903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_104_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_203_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06203_ _01492_ _01478_ _02087_ _02088_ _02089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_118_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07183_ _02650_ _02836_ _02618_ _02837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_195_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06134_ _01953_ _01957_ _02027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_173_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_219_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06065_ _01927_ _01938_ _01944_ _01958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_160_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09824_ soc.rom_encoder_0.request_data_out\[2\] _04743_ _04753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_59_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09755_ _02235_ soc.spi_video_ram_1.write_fifo.fifo_mem\[3\]\[9\] _04697_ _04707_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06967_ _02605_ _02622_ _02627_ _02628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_41_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05918_ _01799_ _01800_ _01796_ _01813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08706_ soc.spi_video_ram_1.fifo_in_address\[6\] _04063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_230_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09686_ soc.rom_encoder_0.request_address\[7\] _04618_ _04659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2106 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_243_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06898_ _02556_ _02560_ _02561_ _00230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_55_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2117 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_214_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2128 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08637_ _04023_ _00506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_15_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2139 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05849_ _01722_ _01738_ _01747_ _01748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_1405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_167_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_230_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_208_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08568_ _02157_ soc.spi_video_ram_1.write_fifo.fifo_mem\[2\]\[18\] _03978_ _03987_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_202_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07519_ _02941_ soc.spi_video_ram_1.write_fifo.fifo_mem\[13\]\[26\] _03167_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_54_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08499_ _03950_ _00441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_22_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_180_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10530_ soc.ram_encoder_0.address\[6\] soc.cpu.AReg.data\[6\] _05227_ _05235_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_196_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xfanout87 soc.cpu.AReg.clk net87 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_50_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_1440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_10_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10461_ soc.cpu.PC.REG.data\[4\] _05183_ _05184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_136_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12200_ _01228_ clknet_leaf_33_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[19\]\[11\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_leaf_280_wb_clk_i clknet_5_4_0_wb_clk_i clknet_leaf_280_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_104_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10392_ _02242_ soc.spi_video_ram_1.write_fifo.fifo_mem\[6\]\[12\] _05135_ _05138_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_124_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12131_ _01159_ clknet_leaf_285_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[6\]\[23\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_174_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_159_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12062_ _01105_ clknet_leaf_108_wb_clk_i soc.rom_loader.current_address\[2\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_111_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11013_ _00079_ clknet_leaf_248_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[16\]\[9\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_89_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_237_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4020 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_133_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_4031 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4042 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4053 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_4064 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_206_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4075 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_219_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4086 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4097 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_233_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_185_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11915_ _00974_ clknet_leaf_121_wb_clk_i soc.cpu.ALU.zx vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_79_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11846_ _00905_ clknet_leaf_166_wb_clk_i soc.rom_encoder_0.request_data_out\[7\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_57_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_221_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1950 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2695 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1961 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1972 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1983 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11777_ _00838_ clknet_leaf_104_wb_clk_i soc.rom_encoder_0.output_buffer\[8\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_207_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1994 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10728_ soc.spi_video_ram_1.write_fifo.fifo_mem\[31\]\[1\] soc.spi_video_ram_1.fifo_in_data\[1\]
+ _05344_ _05346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_147_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10659_ soc.spi_video_ram_1.write_fifo.fifo_mem\[19\]\[28\] soc.spi_video_ram_1.fifo_in_address\[12\]
+ _05277_ _05308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_122_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_1726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12329_ _01357_ clknet_leaf_189_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[8\]\[8\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_138_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_229_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_214_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07870_ _02984_ _03510_ _03513_ _03514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_68_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06821_ _02484_ _02481_ _02497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_110_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09540_ _04558_ _04559_ _00874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_3_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06752_ soc.spi_video_ram_1.write_fifo.fifo_mem\[14\]\[28\] _02353_ _02390_ _02432_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_114_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_225_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05703_ _01588_ _01609_ _01610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
Xclkbuf_leaf_13_wb_clk_i clknet_5_2_0_wb_clk_i clknet_leaf_13_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_92_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09471_ soc.rom_encoder_0.output_buffer\[19\] _04479_ _04516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_77_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_64_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06683_ _02390_ _02391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_92_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_212_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08422_ _03908_ _00406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05634_ _01501_ soc.spi_video_ram_1.output_buffer\[1\] _01543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_225_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_211_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08353_ soc.spi_video_ram_1.write_fifo.fifo_mem\[26\]\[5\] _02401_ _03866_ _03872_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_05565_ soc.spi_video_ram_1.buffer_index\[5\] _01474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_205_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_162_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07304_ _02744_ soc.spi_video_ram_1.write_fifo.fifo_mem\[22\]\[10\] _02954_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_71_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08284_ _03834_ _00342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_138_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05496_ _01409_ _01410_ _01411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_137_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_34_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07235_ soc.spi_video_ram_1.write_fifo.fifo_mem\[8\]\[9\] soc.spi_video_ram_1.write_fifo.fifo_mem\[9\]\[9\]
+ soc.spi_video_ram_1.write_fifo.fifo_mem\[10\]\[9\] soc.spi_video_ram_1.write_fifo.fifo_mem\[11\]\[9\]
+ _02645_ _02614_ _02886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_192_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07166_ _02627_ _02820_ _02821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_117_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_238_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06117_ _01907_ _01975_ _01983_ _01924_ _02010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_69_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_69_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07097_ _02697_ soc.spi_video_ram_1.write_fifo.fifo_mem\[12\]\[3\] _02753_ _02754_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_191_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_117_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06048_ _01939_ _01940_ _01941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_232_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_173_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_219_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09807_ soc.rom_encoder_0.toggled_sram_sck _04737_ _04738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_115_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07999_ _02736_ _03637_ _03638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_189_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09738_ _04698_ _00933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_215_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09669_ soc.cpu.PC.REG.data\[3\] _04646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_231_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_199_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11700_ _00761_ clknet_leaf_198_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[9\]\[2\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_188_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_203_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_180_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11631_ _00009_ clknet_leaf_62_wb_clk_i soc.spi_video_ram_1.current_state\[4\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_145_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_204_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11562_ _00628_ clknet_leaf_293_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[25\]\[27\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_195_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10513_ soc.synch_hack_writeM _05224_ _05225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_11493_ _00559_ clknet_leaf_20_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[24\]\[16\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_11_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xcaravel_hack_soc_110 io_oeb[36] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_10444_ _05170_ _05171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_104_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xcaravel_hack_soc_121 io_out[30] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_104_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_178_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xcaravel_hack_soc_132 la_data_out[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_124_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xcaravel_hack_soc_143 la_data_out[15] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xcaravel_hack_soc_154 la_data_out[26] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_3_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10375_ _02225_ soc.spi_video_ram_1.write_fifo.fifo_mem\[6\]\[4\] _05124_ _05129_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xcaravel_hack_soc_165 la_data_out[38] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xcaravel_hack_soc_176 la_data_out[49] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xcaravel_hack_soc_187 la_data_out[60] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xcaravel_hack_soc_198 wbs_dat_o[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_174_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12114_ _01142_ clknet_leaf_246_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[6\]\[6\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_112_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12045_ net22 clknet_5_31_0_wb_clk_i soc.rom_encoder_0.data_out\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_215_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_78_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_207_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3160 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3171 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_228_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3182 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_244_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11829_ _00888_ clknet_leaf_121_wb_clk_i soc.rom_encoder_0.input_buffer\[3\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1780 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_187_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1791 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_222_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_174_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07020_ _02572_ _02679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_60_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_115_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08971_ soc.spi_video_ram_1.write_fifo.fifo_mem\[22\]\[27\] _02351_ _04177_ _04207_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_233_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_29_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07922_ _02635_ soc.spi_video_ram_1.write_fifo.fifo_mem\[28\]\[21\] _03564_ _02943_
+ _03565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_9_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07853_ _02582_ _03493_ _03496_ _03497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_111_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_42_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06804_ soc.ram_encoder_0.current_state\[2\] _02480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_3
XFILLER_244_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07784_ _03427_ _03428_ _02976_ _03429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_72_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09523_ soc.spi_video_ram_1.initialized soc.video_generator_1.h_count\[1\] _01839_
+ _04547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_37_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06735_ _02423_ _00205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_65_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_213_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09454_ _04500_ _04501_ _04502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06666_ _02165_ soc.spi_video_ram_1.write_fifo.fifo_mem\[12\]\[22\] _02356_ _02381_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XPHY_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_240_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_90_1702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_52_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05617_ _01521_ _01525_ _01526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08405_ soc.spi_video_ram_1.write_fifo.fifo_mem\[27\]\[0\] _02310_ _03899_ _03900_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_40_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_219_wb_clk_i clknet_5_21_0_wb_clk_i clknet_leaf_219_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_09385_ _04430_ _04448_ _00827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_24_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06597_ soc.spi_video_ram_1.fifo_in_address\[4\] _02343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_71_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08336_ _02177_ soc.spi_video_ram_1.write_fifo.fifo_mem\[1\]\[28\] _03830_ _03861_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_90_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05548_ _01451_ _01454_ _01455_ _01457_ _01458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_205_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08267_ soc.ram_encoder_0.request_data_out\[9\] _03789_ _03821_ _03822_ _02510_ _03823_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_193_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05479_ _01381_ _01394_ _00005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_193_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07218_ _02568_ _02869_ _02870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_08198_ _02443_ _02463_ _03767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_14_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07149_ soc.spi_video_ram_1.write_fifo.fifo_mem\[12\]\[5\] soc.spi_video_ram_1.write_fifo.fifo_mem\[13\]\[5\]
+ soc.spi_video_ram_1.write_fifo.fifo_mem\[14\]\[5\] soc.spi_video_ram_1.write_fifo.fifo_mem\[15\]\[5\]
+ _02635_ _02636_ _02804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_195_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10160_ _04995_ _04996_ _01056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_121_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_156_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10091_ soc.ram_encoder_0.request_data_out\[3\] _04930_ _04943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_212_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_210_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_186_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10993_ _00059_ clknet_leaf_76_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[17\]\[18\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_147_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_230_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_208_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_223_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11614_ _00680_ clknet_leaf_239_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[21\]\[21\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_129_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_1398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11545_ _00611_ clknet_leaf_17_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[25\]\[10\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_106_1477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11476_ _00542_ clknet_leaf_270_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[15\]\[28\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_125_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10427_ _05155_ _01181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_48_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_1718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10358_ soc.cpu.ALU.x\[13\] _05109_ _05119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_174_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_151_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10289_ _05071_ _05075_ _05076_ _01105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_238_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_12028_ _01087_ clknet_leaf_74_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[5\]\[16\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_61_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_1426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_226_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_202_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06520_ _02155_ soc.spi_video_ram_1.write_fifo.fifo_mem\[0\]\[17\] _02290_ _02298_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_34_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_222_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06451_ soc.spi_video_ram_1.fifo_in_address\[3\] _02256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xclkbuf_leaf_312_wb_clk_i clknet_5_1_0_wb_clk_i clknet_leaf_312_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_181_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09170_ _02034_ _04325_ _04326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_159_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06382_ _02209_ _00066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08121_ _01836_ soc.video_generator_1.h_count\[6\] _03719_ _03723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_30_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08052_ soc.spi_video_ram_1.write_fifo.fifo_mem\[11\]\[4\] _02399_ _03680_ _03685_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_198_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_200_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07003_ _02589_ _02662_ _02663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_11_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_1_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_192_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_5309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08954_ _04198_ _00648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_131_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07905_ _02656_ _03534_ _03547_ _03548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_4619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08885_ _04161_ _00616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_229_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3907 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3918 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07836_ _03478_ _03479_ _02976_ _03480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_245_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3929 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_211_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_186_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07767_ _02744_ soc.spi_video_ram_1.write_fifo.fifo_mem\[8\]\[15\] _03411_ _03412_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_71_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_1624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09506_ _02260_ soc.cpu.AReg.data\[5\] _04339_ _04538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06718_ soc.spi_video_ram_1.write_fifo.fifo_mem\[14\]\[11\] _02414_ _02412_ _02415_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_129_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07698_ soc.spi_video_ram_1.write_fifo.fifo_mem\[31\]\[24\] _03344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_1661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_246_1679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_198_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_227_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09437_ soc.rom_encoder_0.output_buffer\[12\] _04479_ _04489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_40_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06649_ _02372_ _00170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_53_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_212_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_209_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09368_ soc.spi_video_ram_1.state_sram_clk_counter\[3\] _04437_ _04433_ _04440_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_21_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_138_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08319_ _03852_ _00359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_138_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09299_ _02225_ soc.spi_video_ram_1.write_fifo.fifo_mem\[4\]\[4\] _04395_ _04400_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_103_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11330_ _00396_ clknet_leaf_297_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[26\]\[27\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_158_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_192_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11261_ _00327_ clknet_leaf_150_wb_clk_i soc.ram_encoder_0.output_buffer\[7\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_108_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10212_ _02221_ soc.spi_video_ram_1.write_fifo.fifo_mem\[5\]\[2\] _05030_ _05033_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_6500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_180_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11192_ _00258_ clknet_leaf_137_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[11\]\[2\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_161_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_6511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_122_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_175_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10143_ soc.ram_encoder_0.request_data_out\[15\] _04929_ _04983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_122_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_171_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_216_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5810 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5821 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5832 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5843 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10074_ _02484_ _02490_ _04929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_94_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5854 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5865 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_47_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_5876 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_130_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5887 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_208_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5898 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_130_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_235_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10976_ _00042_ clknet_leaf_217_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[17\]\[1\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_204_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_231_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_188_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_157_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_129_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11528_ _00594_ clknet_leaf_240_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[23\]\[22\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_7_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11459_ _00525_ clknet_leaf_33_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[15\]\[11\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_113_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_1545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_98_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_193_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_239_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05951_ soc.video_generator_1.h_count\[5\] _01843_ _01844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_23_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08670_ soc.spi_video_ram_1.write_fifo.fifo_mem\[15\]\[8\] _02407_ _04032_ _04041_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_05882_ _01654_ _01769_ _01778_ _01779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
XFILLER_227_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_213_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07621_ _02752_ soc.spi_video_ram_1.write_fifo.fifo_mem\[8\]\[25\] _03267_ _03268_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_94_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07552_ soc.spi_video_ram_1.write_fifo.fifo_mem\[31\]\[13\] _03199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_78_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06503_ _02138_ soc.spi_video_ram_1.write_fifo.fifo_mem\[0\]\[9\] _02279_ _02289_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_35_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07483_ soc.spi_video_ram_1.write_fifo.fifo_mem\[7\]\[12\] _03131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_165_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09222_ _04054_ _04339_ _04357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06434_ soc.spi_video_ram_1.write_fifo.fifo_mem\[16\]\[13\] _02244_ _02238_ _02245_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_107_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_210_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_206_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_1390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09153_ _01866_ _01959_ _03712_ _04313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_06365_ _02155_ soc.spi_video_ram_1.write_fifo.fifo_mem\[17\]\[17\] _02193_ _02201_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_08104_ _01836_ _01968_ _01993_ _03711_ _03712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_120_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09084_ _04272_ _00704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_175_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06296_ soc.spi_video_ram_1.fifo_in_address\[3\] _02159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_174_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08035_ _02685_ _03672_ _02720_ _03673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_163_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_190_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_162_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_115_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5106 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09986_ soc.ram_step2_read_request soc.ram_step1_write_request _02053_ _04875_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_5117 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5128 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5139 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_233_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08937_ soc.spi_video_ram_1.write_fifo.fifo_mem\[22\]\[10\] _02411_ _04189_ _04190_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_4416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_170_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3704 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08868_ _04152_ _00608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3715 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3726 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3737 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_217_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3748 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_234_wb_clk_i clknet_5_16_0_wb_clk_i clknet_leaf_234_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_2_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07819_ soc.spi_video_ram_1.write_fifo.fifo_mem\[15\]\[23\] _03464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_3759 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08799_ _04115_ _00576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_72_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_244_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10830_ _02256_ soc.spi_video_ram_1.write_fifo.fifo_mem\[7\]\[19\] _05389_ _05401_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_25_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10761_ soc.spi_video_ram_1.write_fifo.fifo_mem\[31\]\[16\] soc.spi_video_ram_1.fifo_in_address\[0\]
+ _05355_ _05364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_213_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_224_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10692_ soc.spi_video_ram_1.fifo_in_data\[13\] _05325_ _05327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_125_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_199_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_197_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_240_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_181_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_225_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_194_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_193_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11313_ _00379_ clknet_leaf_17_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[26\]\[10\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12293_ _01321_ clknet_leaf_80_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[7\]\[17\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_154_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11244_ _00310_ clknet_leaf_3_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[10\]\[15\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_84_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_171_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_175_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11175_ _00241_ clknet_leaf_56_wb_clk_i soc.spi_video_ram_1.output_buffer\[15\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_6330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_68_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_6341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_1420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10126_ _04952_ _04970_ _01048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_6374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_114_1510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_5640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_95_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_23_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10057_ _04914_ _01036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_76_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_5684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_209_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_212_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5695 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4950 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4961 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4972 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4983 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_1549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_4994 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_149_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10959_ _00025_ clknet_leaf_40_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[18\]\[13\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_143_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_176_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_223_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06150_ _01967_ _02005_ _02043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xclkbuf_leaf_38_wb_clk_i clknet_5_3_0_wb_clk_i clknet_leaf_38_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_160_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_185_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06081_ _01925_ _01973_ _01974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_172_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_172_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_236_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09840_ soc.rom_encoder_0.request_data_out\[5\] _04743_ _04766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_98_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_58_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09771_ _04715_ _00949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_6_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06983_ _02642_ _02643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_246_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_85_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_230_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08722_ soc.spi_video_ram_1.write_fifo.fifo_mem\[15\]\[28\] _02353_ _04043_ _04073_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_05934_ _01807_ _01810_ _01828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_26_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_05865_ _01754_ _01756_ _01762_ _01763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_08653_ _04031_ _04032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_82_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_226_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07604_ _02575_ soc.spi_video_ram_1.write_fifo.fifo_mem\[28\]\[25\] _03250_ _02943_
+ _03251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_96_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05796_ _01682_ _01695_ _01697_ _01698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08584_ _02173_ soc.spi_video_ram_1.write_fifo.fifo_mem\[2\]\[26\] _03966_ _03995_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_81_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_242_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07535_ _03173_ _03182_ _02567_ _03183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_228_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xclkbuf_2_2_0_wb_clk_i clknet_0_wb_clk_i clknet_2_2_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_07466_ _02607_ soc.spi_video_ram_1.write_fifo.fifo_mem\[20\]\[12\] _03113_ _02943_
+ _03114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_161_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_179_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06417_ soc.spi_video_ram_1.fifo_in_data\[8\] _02233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_09205_ _00011_ _01699_ _04348_ _00749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_241_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07397_ _03041_ _03042_ _03045_ _02570_ _03046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_72_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_176_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06348_ _02138_ soc.spi_video_ram_1.write_fifo.fifo_mem\[17\]\[9\] _02182_ _02192_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_09136_ soc.spi_video_ram_1.state_counter\[5\] _04300_ _04302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_176_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_202_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09067_ _04263_ _00696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06279_ _02147_ soc.spi_video_ram_1.write_fifo.fifo_mem\[18\]\[13\] _02141_ _02148_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_151_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_191_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08018_ _03596_ _03655_ _03656_ _00254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_239_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_176_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09969_ soc.ram_encoder_0.input_buffer\[7\] _04863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_4202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_213_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11931_ _00990_ clknet_leaf_164_wb_clk_i soc.ram_encoder_0.input_bits_left\[2\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_4279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2800 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_175_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2811 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2822 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2833 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11862_ _00921_ clknet_leaf_109_wb_clk_i soc.rom_encoder_0.request_address\[7\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2844 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2855 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2866 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_207_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10813_ _05391_ _01315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2877 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2888 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2899 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11793_ _00854_ clknet_leaf_130_wb_clk_i soc.spi_video_ram_1.buffer_index\[4\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_232_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10744_ soc.spi_video_ram_1.write_fifo.fifo_mem\[31\]\[9\] soc.spi_video_ram_1.fifo_in_data\[9\]
+ _05344_ _05354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_186_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_185_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10675_ _02229_ soc.spi_video_ram_1.write_fifo.fifo_mem\[29\]\[6\] _05310_ _05317_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_139_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_220_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12345_ _01373_ clknet_leaf_306_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[8\]\[24\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_103_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12276_ _01304_ clknet_leaf_213_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[7\]\[0\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_107_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_194_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_155_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11227_ _00293_ clknet_leaf_85_wb_clk_i soc.video_generator_1.h_count\[8\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_136_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_218_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6160 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11158_ _00224_ net84 soc.cpu.AReg.data\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_leaf_156_wb_clk_i clknet_5_30_0_wb_clk_i clknet_leaf_156_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_150_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6171 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6182 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_23_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10109_ soc.ram_data_out\[6\] _04927_ _04957_ _04958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_231_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11089_ _00155_ clknet_leaf_41_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[13\]\[27\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_5470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_7_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_236_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4780 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_110_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_208_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4791 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05650_ soc.cpu.ALU.zx _01558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_36_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_224_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_210_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05581_ soc.spi_video_ram_1.output_buffer\[11\] soc.spi_video_ram_1.output_buffer\[10\]
+ _01461_ _01490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_229_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_177_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07320_ _00003_ _02970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_32_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07251_ _02572_ _02902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_220_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06202_ _01492_ _01481_ _02088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07182_ soc.spi_video_ram_1.write_fifo.fifo_mem\[4\]\[6\] soc.spi_video_ram_1.write_fifo.fifo_mem\[5\]\[6\]
+ soc.spi_video_ram_1.write_fifo.fifo_mem\[6\]\[6\] soc.spi_video_ram_1.write_fifo.fifo_mem\[7\]\[6\]
+ _02613_ _02652_ _02836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_191_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_157_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_203_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06133_ _02003_ _02023_ _02025_ _02026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_173_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06064_ _01954_ _01955_ _01956_ _01957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_67_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09823_ _01395_ _04752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_134_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_246_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_150_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09754_ _04706_ _00941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_86_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06966_ _01411_ _02626_ _02627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_228_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08705_ _03541_ _04046_ _04062_ _00535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_05917_ _01805_ _01798_ _01811_ _01812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_09685_ _04639_ soc.rom_loader.current_address\[7\] _04657_ _04658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06897_ soc.ram_encoder_0.output_buffer\[3\] _02558_ _02561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_54_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2107 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2118 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2129 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_227_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08636_ _02163_ soc.spi_video_ram_1.write_fifo.fifo_mem\[30\]\[21\] _03999_ _04023_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_76_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05848_ _01746_ _01747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_1406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_243_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08567_ _03986_ _00473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_120_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_214_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05779_ _01594_ _01680_ _01681_ _01590_ soc.cpu.PC.in\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_23_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07518_ soc.spi_video_ram_1.write_fifo.fifo_mem\[8\]\[26\] soc.spi_video_ram_1.write_fifo.fifo_mem\[9\]\[26\]
+ soc.spi_video_ram_1.write_fifo.fifo_mem\[10\]\[26\] soc.spi_video_ram_1.write_fifo.fifo_mem\[11\]\[26\]
+ _02783_ _02690_ _03166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_126_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_167_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08498_ _02149_ soc.spi_video_ram_1.write_fifo.fifo_mem\[28\]\[14\] _03945_ _03950_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_126_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_208_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_221_1722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout88 net89 net88 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_07449_ _02696_ soc.spi_video_ram_1.write_fifo.fifo_mem\[28\]\[27\] _03097_ _03098_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_17_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_210_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10460_ _04646_ _05180_ _05183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_149_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09119_ soc.spi_video_ram_1.current_state\[2\] _04290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_10391_ _05137_ _01147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_237_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12130_ _01158_ clknet_leaf_269_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[6\]\[22\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_150_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12061_ _01104_ clknet_leaf_107_wb_clk_i soc.rom_loader.current_address\[1\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_46_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11012_ _00078_ clknet_leaf_218_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[16\]\[8\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_46_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_1286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4010 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4021 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4032 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4043 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4054 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4065 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_218_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4076 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4087 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4098 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11914_ _00973_ clknet_leaf_128_wb_clk_i soc.cpu.ALU.nx vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_59_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_206_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11845_ _00904_ clknet_leaf_169_wb_clk_i soc.rom_encoder_0.request_data_out\[6\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1940 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_220_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1951 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_233_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2696 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1962 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1973 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11776_ _00837_ clknet_leaf_93_wb_clk_i soc.rom_encoder_0.output_buffer\[7\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_14_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1984 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1995 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_198_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10727_ _05345_ _01275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_202_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10658_ _05307_ _01244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_70_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10589_ _05266_ _05268_ _05269_ _01213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_170_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12328_ _01356_ clknet_leaf_193_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[8\]\[7\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_170_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12259_ _01287_ clknet_leaf_311_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[31\]\[12\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_68_1492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_1462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_69_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_190_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_151_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06820_ soc.ram_encoder_0.output_bits_left\[3\] soc.ram_encoder_0.output_bits_left\[2\]
+ _02496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_99_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06751_ _02431_ _00213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_243_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_237_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_92_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_184_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05702_ _01562_ _01597_ _01607_ _01609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_37_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_209_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09470_ soc.rom_encoder_0.output_buffer\[15\] _02455_ _04514_ _02461_ _04515_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_52_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06682_ _02389_ _02390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_227_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_225_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_221_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08421_ soc.spi_video_ram_1.write_fifo.fifo_mem\[27\]\[8\] _02407_ _03899_ _03908_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_145_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05633_ _01541_ _01542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_196_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_205_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xclkbuf_leaf_53_wb_clk_i clknet_5_13_0_wb_clk_i clknet_leaf_53_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_05564_ _01468_ _01471_ _01472_ _01473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_08352_ _03871_ _00373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_149_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07303_ _02758_ _02948_ _02951_ _02952_ _02953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_138_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08283_ _02124_ soc.spi_video_ram_1.write_fifo.fifo_mem\[1\]\[2\] _03831_ _03834_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_05495_ soc.spi_video_ram_1.current_state\[1\] soc.spi_video_ram_1.current_state\[4\]
+ _01410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_20_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07234_ _02650_ _02884_ _02885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_146_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07165_ _02606_ _02810_ _02819_ _02820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_30_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_118_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_246_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06116_ _02004_ _02008_ _02009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_118_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_173_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07096_ _02752_ soc.spi_video_ram_1.write_fifo.fifo_mem\[13\]\[3\] _02753_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_246_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06047_ _01853_ _01850_ _01940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_82_1423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09806_ _04736_ _02463_ _04566_ _04571_ _04737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_86_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07998_ soc.spi_video_ram_1.write_fifo.fifo_mem\[8\]\[17\] soc.spi_video_ram_1.write_fifo.fifo_mem\[9\]\[17\]
+ soc.spi_video_ram_1.write_fifo.fifo_mem\[10\]\[17\] soc.spi_video_ram_1.write_fifo.fifo_mem\[11\]\[17\]
+ _02701_ _02737_ _03637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_235_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_214_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09737_ _02213_ soc.spi_video_ram_1.write_fifo.fifo_mem\[3\]\[0\] _04697_ _04698_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_21_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06949_ soc.spi_video_ram_1.write_fifo.fifo_mem\[24\]\[0\] soc.spi_video_ram_1.write_fifo.fifo_mem\[25\]\[0\]
+ soc.spi_video_ram_1.write_fifo.fifo_mem\[26\]\[0\] soc.spi_video_ram_1.write_fifo.fifo_mem\[27\]\[0\]
+ _02607_ _02578_ _02610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_55_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09668_ _04645_ _00916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_27_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08619_ _04014_ _00497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_82_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09599_ _01380_ _04601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_202_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_215_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11630_ _00008_ clknet_leaf_64_wb_clk_i soc.spi_video_ram_1.current_state\[3\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_54_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11561_ _00627_ clknet_leaf_292_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[25\]\[26\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_138_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_126_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10512_ _05218_ soc.hack_clk_strobe _05223_ _05224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_13_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11492_ _00558_ clknet_leaf_313_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[24\]\[15\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_7_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_196_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xcaravel_hack_soc_100 io_oeb[9] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xcaravel_hack_soc_111 io_oeb[37] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_10443_ soc.cpu.DMuxJMP.sel\[2\] _02539_ _05165_ _05169_ _01552_ _05170_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai221_4
XFILLER_6_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xcaravel_hack_soc_122 io_out[31] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_13_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_100_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xcaravel_hack_soc_133 la_data_out[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_137_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xcaravel_hack_soc_144 la_data_out[16] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_174_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xcaravel_hack_soc_155 la_data_out[28] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xcaravel_hack_soc_166 la_data_out[39] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_174_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10374_ _05128_ _01139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xcaravel_hack_soc_177 la_data_out[50] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_151_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xcaravel_hack_soc_188 la_data_out[61] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_12113_ _01141_ clknet_leaf_245_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[6\]\[5\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xcaravel_hack_soc_199 wbs_dat_o[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_65_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12044_ net21 clknet_leaf_87_wb_clk_i soc.rom_encoder_0.data_out\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_46_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_211_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_232_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_225_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_219_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_185_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3150 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3161 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3172 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3183 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_207_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_1349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_209_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_221_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11828_ _00887_ clknet_leaf_124_wb_clk_i soc.rom_encoder_0.input_buffer\[2\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_187_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1781 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1792 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11759_ _00820_ clknet_leaf_71_wb_clk_i soc.spi_video_ram_1.state_sram_clk_counter\[2\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_14_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_220_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_100_wb_clk_i clknet_5_14_0_wb_clk_i clknet_leaf_100_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_08970_ _04206_ _00656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_130_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07921_ _02931_ _03563_ _03564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_116_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07852_ _02752_ soc.spi_video_ram_1.write_fifo.fifo_mem\[28\]\[22\] _03495_ _02927_
+ _03496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_60_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_217_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06803_ soc.ram_encoder_0.output_bits_left\[4\] _02478_ _02479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_84_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput1 io_in[10] net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_211_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07783_ _02926_ soc.spi_video_ram_1.write_fifo.fifo_mem\[16\]\[23\] _03428_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_186_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09522_ _01994_ soc.video_generator_1.h_count\[4\] soc.video_generator_1.h_count\[7\]
+ _04546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_06734_ soc.spi_video_ram_1.write_fifo.fifo_mem\[14\]\[19\] _02341_ _02412_ _02423_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_83_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09453_ _02458_ _03766_ soc.rom_encoder_0.output_buffer\[12\] _04501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06665_ _02380_ _00178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_64_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_164_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_08404_ _03898_ _03899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_197_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05616_ _01471_ _01522_ _01523_ _01524_ _01525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_75_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09384_ _04448_ _04450_ _00826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06596_ _02342_ _00147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_75_1282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08335_ _03860_ _00367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_244_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05547_ net87 soc.hack_clk_strobe soc.cpu.AReg.data\[14\] _01456_ _01457_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_36_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_137_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08266_ soc.ram_encoder_0.output_buffer\[13\] _03817_ _03822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_05478_ soc.spi_video_ram_1.current_state\[0\] _01393_ _01394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_193_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_192_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xclkbuf_leaf_259_wb_clk_i clknet_5_18_0_wb_clk_i clknet_leaf_259_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_197_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07217_ _02862_ _02864_ _02866_ _02868_ _02869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_118_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08197_ _02445_ _03765_ _03766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_106_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_238_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_119_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_84_1507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07148_ _02583_ _02802_ _02803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_161_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_156_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07079_ _02643_ _02736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_161_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10090_ _04787_ _04942_ _01040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_207_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10992_ _00058_ clknet_leaf_79_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[17\]\[17\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_186_1753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_231_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_147_1726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_167_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_203_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_187_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11613_ _00679_ clknet_leaf_50_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[21\]\[20\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_204_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11544_ _00610_ clknet_leaf_257_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[25\]\[9\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_184_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_183_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11475_ _00541_ clknet_leaf_42_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[15\]\[27\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_125_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10426_ _01378_ _05016_ _05155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_67_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_152_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10357_ _01803_ _05104_ _05118_ _01132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_139_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_174_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_215_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10288_ soc.rom_loader.current_address\[2\] soc.rom_loader.current_address\[1\] _05069_
+ _05076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_111_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_12027_ _01086_ clknet_leaf_312_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[5\]\[15\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_78_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_65_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_228_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06450_ _02255_ _00088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_181_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_107_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_241_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_222_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_163_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06381_ _02171_ soc.spi_video_ram_1.write_fifo.fifo_mem\[17\]\[25\] _02181_ _02209_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_37_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_241_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08120_ _01836_ _03719_ soc.video_generator_1.h_count\[6\] _03722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_119_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_174_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_1753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08051_ _03684_ _00259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_239_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07002_ soc.spi_video_ram_1.write_fifo.fifo_mem\[16\]\[1\] soc.spi_video_ram_1.write_fifo.fifo_mem\[17\]\[1\]
+ soc.spi_video_ram_1.write_fifo.fifo_mem\[18\]\[1\] soc.spi_video_ram_1.write_fifo.fifo_mem\[19\]\[1\]
+ _02645_ _02614_ _02662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_115_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08953_ soc.spi_video_ram_1.write_fifo.fifo_mem\[22\]\[18\] _02339_ _04189_ _04198_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_170_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07904_ _02831_ _03540_ _03546_ _03547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_97_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08884_ soc.spi_video_ram_1.write_fifo.fifo_mem\[25\]\[15\] _04054_ _04155_ _04161_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_3908 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07835_ _03021_ soc.spi_video_ram_1.write_fifo.fifo_mem\[16\]\[22\] _03479_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_116_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3919 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_244_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_42_1281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_186_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07766_ _03139_ _03410_ _03411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_65_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09505_ _04537_ _00861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_53_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06717_ soc.spi_video_ram_1.fifo_in_data\[11\] _02414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_213_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_246_1647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07697_ soc.spi_video_ram_1.write_fifo.fifo_mem\[24\]\[24\] soc.spi_video_ram_1.write_fifo.fifo_mem\[25\]\[24\]
+ soc.spi_video_ram_1.write_fifo.fifo_mem\[26\]\[24\] soc.spi_video_ram_1.write_fifo.fifo_mem\[27\]\[24\]
+ _02902_ _02576_ _03343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_52_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_240_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09436_ soc.rom_encoder_0.request_address\[11\] _02520_ _04460_ soc.rom_encoder_0.output_buffer\[8\]
+ _04487_ _04488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XPHY_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_06648_ _02147_ soc.spi_video_ram_1.write_fifo.fifo_mem\[12\]\[13\] _02368_ _02372_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_52_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_80_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_201_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09367_ soc.spi_video_ram_1.state_sram_clk_counter\[3\] _04437_ _04439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_234_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_166_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06579_ soc.spi_video_ram_1.write_fifo.fifo_mem\[13\]\[13\] _02244_ _02328_ _02332_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_205_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08318_ _02159_ soc.spi_video_ram_1.write_fifo.fifo_mem\[1\]\[19\] _03842_ _03852_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_166_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09298_ _04399_ _00791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_90_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_193_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_165_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08249_ soc.ram_encoder_0.request_address\[13\] _02505_ _03808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_14_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_88_1451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11260_ _00326_ clknet_leaf_150_wb_clk_i soc.ram_encoder_0.output_buffer\[6\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_10_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_107_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10211_ _05032_ _01072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_218_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11191_ _00257_ clknet_leaf_190_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[11\]\[1\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_6501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_234_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10142_ _04952_ _04982_ _01052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_6534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5800 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5811 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5822 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5833 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10073_ _04926_ _04928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_121_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_212_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_6589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5844 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5855 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_236_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5866 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_134_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5877 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5888 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5899 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10975_ _00041_ clknet_5_23_0_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[17\]\[0\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_189_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_245_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_223_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_156_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11527_ _00593_ clknet_leaf_240_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[23\]\[21\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_106_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11458_ _00524_ clknet_leaf_15_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[15\]\[10\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_67_1513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10409_ _05146_ _01156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_139_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_3_4_0_wb_clk_i clknet_2_2_0_wb_clk_i clknet_3_4_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_113_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11389_ _00455_ clknet_leaf_303_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[28\]\[28\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_113_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05950_ soc.video_generator_1.h_count\[3\] soc.video_generator_1.h_count\[4\] _01842_
+ _01843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_05881_ _01775_ _01777_ _01778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_226_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07620_ _02763_ _03266_ _03267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_19_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_242_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07551_ soc.spi_video_ram_1.write_fifo.fifo_mem\[24\]\[13\] soc.spi_video_ram_1.write_fifo.fifo_mem\[25\]\[13\]
+ soc.spi_video_ram_1.write_fifo.fifo_mem\[26\]\[13\] soc.spi_video_ram_1.write_fifo.fifo_mem\[27\]\[13\]
+ _03139_ _02908_ _03198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_74_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06502_ _02288_ _00107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_222_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07482_ _02613_ soc.spi_video_ram_1.write_fifo.fifo_mem\[4\]\[12\] _03129_ _02943_
+ _03130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_22_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09221_ _04341_ _01834_ _04356_ _00757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06433_ soc.spi_video_ram_1.fifo_in_data\[13\] _02244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_22_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09152_ _04294_ _04312_ _00732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06364_ _02200_ _00057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_202_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_148_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_124_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08103_ soc.video_generator_1.h_count\[4\] soc.video_generator_1.h_count\[7\] soc.video_generator_1.h_count\[6\]
+ _03711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_147_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09083_ _02240_ soc.spi_video_ram_1.write_fifo.fifo_mem\[20\]\[11\] _04270_ _04272_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06295_ _02158_ _00030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_198_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_200_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08034_ soc.spi_video_ram_1.write_fifo.fifo_mem\[20\]\[16\] soc.spi_video_ram_1.write_fifo.fifo_mem\[21\]\[16\]
+ soc.spi_video_ram_1.write_fifo.fifo_mem\[22\]\[16\] soc.spi_video_ram_1.write_fifo.fifo_mem\[23\]\[16\]
+ _02717_ _02682_ _03672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_176_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_137_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_192_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_235_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09985_ _02484_ _02498_ _04874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_103_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_5107 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5118 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_130_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5129 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08936_ _04176_ _04189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_88_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_213_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_229_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_218_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08867_ soc.spi_video_ram_1.write_fifo.fifo_mem\[25\]\[7\] _02405_ _04144_ _04152_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_3705 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3716 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3727 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3738 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07818_ _03458_ _03459_ _03462_ _02691_ _02929_ _03463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XTAP_3749 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08798_ _02128_ soc.spi_video_ram_1.write_fifo.fifo_mem\[23\]\[4\] _04110_ _04115_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_84_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_8_wb_clk_i clknet_5_2_0_wb_clk_i clknet_leaf_8_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_07749_ _02893_ _03393_ _03394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_60_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_26_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_241_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_198_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10760_ _03393_ _05358_ _05363_ _01290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_242_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_274_wb_clk_i clknet_5_6_0_wb_clk_i clknet_leaf_274_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_1481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_246_1488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09419_ soc.rom_encoder_0.request_address\[7\] _02520_ _04460_ soc.rom_encoder_0.output_buffer\[4\]
+ _04474_ _04475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_10691_ _03118_ _05324_ _05326_ _01258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xclkbuf_leaf_203_wb_clk_i clknet_5_22_0_wb_clk_i clknet_leaf_203_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_90_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_200_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_1404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_126_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_218_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_11312_ _00378_ clknet_leaf_259_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[26\]\[9\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_5_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12292_ _01320_ clknet_leaf_75_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[7\]\[16\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_154_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11243_ _00309_ clknet_leaf_6_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[10\]\[14\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_122_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_190_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11174_ _00240_ clknet_5_24_0_wb_clk_i soc.spi_video_ram_1.output_buffer\[16\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_6331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10125_ soc.ram_data_out\[10\] _04928_ _04969_ _04970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_6364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_1465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10056_ soc.ram_encoder_0.request_address\[14\] soc.ram_encoder_0.address\[14\] _04879_
+ _04914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_5674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_208_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4940 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_1498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_5696 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4951 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4962 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_4973 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_114_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_235_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_224_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_188_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4984 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4995 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_169_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_204_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10958_ _00024_ clknet_leaf_2_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[18\]\[12\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_182_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_231_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_188_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_108_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_189_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10889_ soc.spi_video_ram_1.write_fifo.fifo_mem\[8\]\[1\] soc.spi_video_ram_1.fifo_in_data\[1\]
+ _05431_ _05433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XPHY_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_157_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_31_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_201_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06080_ soc.display_clks_before_active\[0\] soc.video_generator_1.h_count\[2\] _01903_
+ _01967_ _01973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or4_1
XFILLER_176_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_208_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_78_wb_clk_i clknet_5_8_0_wb_clk_i clknet_leaf_78_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_98_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_193_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_217_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09770_ _02250_ soc.spi_video_ram_1.write_fifo.fifo_mem\[3\]\[16\] _04708_ _04715_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06982_ _00002_ _02642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_67_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08721_ _04072_ _00541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05933_ _01816_ _01815_ _01826_ _01827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XTAP_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_227_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08652_ soc.spi_video_ram_1.write_fifo.write_pointer\[4\] _01449_ _04031_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_05864_ _01758_ _01761_ _01762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_66_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07603_ _03054_ _03249_ _03250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08583_ _03994_ _00481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05795_ _01586_ _01696_ _01697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_82_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07534_ _02984_ _03174_ _03181_ _02601_ _03182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_23_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_223_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_243_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07465_ _03054_ _03112_ _03113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_210_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_206_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09204_ soc.spi_video_ram_1.fifo_in_data\[6\] _04346_ _04348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06416_ _02232_ _00077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_22_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07396_ _03043_ _03044_ _02958_ _03045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_52_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09135_ _04294_ _04300_ _04301_ _00726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_136_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06347_ _02191_ _00049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_104_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09066_ _02223_ soc.spi_video_ram_1.write_fifo.fifo_mem\[20\]\[3\] _04259_ _04263_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06278_ soc.spi_video_ram_1.fifo_in_data\[13\] _02147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_120_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_190_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_159_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08017_ soc.spi_video_ram_1.output_buffer\[2\] _02675_ _03656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_102_1492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_131_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09968_ _04861_ _04848_ _04862_ _00999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_76_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08919_ _04180_ _00631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_170_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09899_ _02454_ _04810_ _04811_ _00981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_4236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_4247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11930_ _00989_ clknet_leaf_160_wb_clk_i soc.ram_encoder_0.toggled_sram_sck vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_2
XTAP_4258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_217_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_206_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2801 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2812 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2823 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11861_ _00920_ clknet_leaf_105_wb_clk_i soc.rom_encoder_0.request_address\[6\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2834 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_168_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2845 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2856 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10812_ _02240_ soc.spi_video_ram_1.write_fifo.fifo_mem\[7\]\[11\] _05389_ _05391_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_2867 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2878 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11792_ _00853_ clknet_leaf_130_wb_clk_i soc.spi_video_ram_1.buffer_index\[3\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_26_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2889 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_213_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_183_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_159_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10743_ _05353_ _01283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_159_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_201_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10674_ _05316_ _01251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_139_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_185_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12344_ _01372_ clknet_leaf_238_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[8\]\[23\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_99_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_12275_ _01303_ clknet_leaf_303_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[31\]\[28\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_120_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11226_ _00292_ clknet_leaf_86_wb_clk_i soc.video_generator_1.h_count\[7\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_136_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_6150 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11157_ _00223_ clknet_leaf_95_wb_clk_i soc.rom_encoder_0.output_bits_left\[2\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_150_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6161 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_155_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6172 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6183 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10108_ _04853_ _04947_ _04948_ _04956_ _04957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_110_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11088_ _00154_ clknet_leaf_279_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[13\]\[26\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_209_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10039_ _04905_ _01027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xclkbuf_leaf_196_wb_clk_i clknet_5_25_0_wb_clk_i clknet_leaf_196_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_4770 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4781 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4792 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_125_wb_clk_i clknet_5_12_0_wb_clk_i clknet_leaf_125_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_64_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_205_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05580_ _01478_ _01482_ _01483_ _01484_ _01486_ _01488_ _01489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_189_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_5_25_0_wb_clk_i clknet_4_12_0_wb_clk_i clknet_5_25_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_177_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_20_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_182_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07250_ _02900_ _02901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_83_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_158_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_223_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_1350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06201_ _01470_ _01494_ _02087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_125_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07181_ _02589_ _02834_ _02835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_160_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_219_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06132_ _01954_ _02024_ _02025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_117_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_172_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06063_ _01848_ _01890_ _01916_ _01918_ _01919_ _01956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_86_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_105_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_236_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_63_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09822_ _01396_ _04751_ _00964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_58_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_214_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_80_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09753_ _02233_ soc.spi_video_ram_1.write_fifo.fifo_mem\[3\]\[8\] _04697_ _04706_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_230_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06965_ _02623_ _02625_ _02626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_171_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08704_ _04061_ _04048_ _04062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05916_ _01807_ _01810_ _01811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_27_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09684_ _04639_ _04656_ _04657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06896_ soc.ram_encoder_0.request_address\[2\] _02506_ _02560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2108 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2119 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08635_ _04022_ _00505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05847_ _01744_ _01745_ _01746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_55_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_242_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08566_ _02155_ soc.spi_video_ram_1.write_fifo.fifo_mem\[2\]\[17\] _03978_ _03986_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_05778_ _01553_ soc.cpu.AReg.data\[5\] _01681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07517_ _03155_ _03164_ _03165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_126_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08497_ _03949_ _00440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_50_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_211_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_168_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07448_ _02612_ soc.spi_video_ram_1.write_fifo.fifo_mem\[29\]\[27\] _03097_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_74_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_156_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout89 net90 net89 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_109_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07379_ _03021_ soc.spi_video_ram_1.write_fifo.fifo_mem\[23\]\[11\] _02614_ _03028_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_136_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_202_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09118_ _04289_ _00721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_129_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10390_ _02240_ soc.spi_video_ram_1.write_fifo.fifo_mem\[6\]\[11\] _05135_ _05137_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_139_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09049_ _04243_ _04250_ _04251_ _00690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_191_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12060_ _01103_ clknet_leaf_107_wb_clk_i soc.rom_loader.current_address\[0\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_104_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11011_ _00077_ clknet_leaf_187_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[16\]\[7\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_150_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_4000 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4011 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_77_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4022 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_4033 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_213_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4044 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4055 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4066 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4077 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11913_ _00972_ clknet_5_26_0_wb_clk_i soc.cpu.ALU.zy vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_4088 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4099 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_234_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11844_ _00903_ clknet_leaf_95_wb_clk_i soc.rom_encoder_0.request_data_out\[5\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1930 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1941 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1952 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2697 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1963 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11775_ _00836_ clknet_leaf_107_wb_clk_i soc.rom_encoder_0.output_buffer\[6\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_226_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1974 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1985 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1996 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10726_ soc.spi_video_ram_1.write_fifo.fifo_mem\[31\]\[0\] soc.spi_video_ram_1.fifo_in_data\[0\]
+ _05344_ _05345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_179_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10657_ soc.spi_video_ram_1.write_fifo.fifo_mem\[19\]\[27\] soc.spi_video_ram_1.fifo_in_address\[11\]
+ _05277_ _05307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_220_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_167_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10588_ soc.gpio_i_stored\[0\] _05268_ _02053_ _05269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_103_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_154_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12327_ _01355_ clknet_leaf_205_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[8\]\[6\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_157_1728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_126_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12258_ _01286_ clknet_leaf_37_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[31\]\[11\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_218_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11209_ _00275_ clknet_leaf_30_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[11\]\[19\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_68_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12189_ _01217_ clknet_leaf_189_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[19\]\[0\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_96_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_231_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xclkbuf_leaf_306_wb_clk_i clknet_5_3_0_wb_clk_i clknet_leaf_306_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_7_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06750_ soc.spi_video_ram_1.write_fifo.fifo_mem\[14\]\[27\] _02351_ _02390_ _02431_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_83_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_236_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05701_ _01561_ _01607_ _01608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_06681_ _02388_ _02314_ _02389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_63_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_110_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08420_ _03907_ _00405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_224_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05632_ _01501_ _01539_ _01540_ _01470_ _01541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_91_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_244_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_229_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08351_ soc.spi_video_ram_1.write_fifo.fifo_mem\[26\]\[4\] _02399_ _03866_ _03871_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_05563_ _01461_ soc.spi_video_ram_1.buffer_index\[1\] _01470_ _01472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_166_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_1317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07302_ _02581_ _02952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_08282_ _03833_ _00341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05494_ soc.spi_video_ram_1.current_state\[3\] _01409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_220_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07233_ soc.spi_video_ram_1.write_fifo.fifo_mem\[12\]\[9\] soc.spi_video_ram_1.write_fifo.fifo_mem\[13\]\[9\]
+ soc.spi_video_ram_1.write_fifo.fifo_mem\[14\]\[9\] soc.spi_video_ram_1.write_fifo.fifo_mem\[15\]\[9\]
+ _02645_ _02614_ _02884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
Xclkbuf_leaf_93_wb_clk_i clknet_5_14_0_wb_clk_i clknet_leaf_93_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_149_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_203_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_22_wb_clk_i clknet_5_8_0_wb_clk_i clknet_leaf_22_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_07164_ _02812_ _02814_ _02816_ _02818_ _02620_ _02819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_101_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06115_ _01986_ _02006_ _02007_ _01977_ _02008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_173_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07095_ _02574_ _02752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_145_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06046_ soc.video_generator_1.v_count\[5\] _01939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_132_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_1446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09805_ _02445_ _04736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_60_1722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07997_ _03596_ _03635_ _03636_ _00253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_228_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_46_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09736_ _04696_ _04697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_06948_ _02596_ _02608_ _02609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_210_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09667_ _04644_ soc.rom_encoder_0.request_address\[2\] _04632_ _04645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_227_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06879_ soc.rom_encoder_0.output_buffer\[2\] _02542_ _02543_ soc.rom_encoder_0.request_address\[1\]
+ _02546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_216_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08618_ _02145_ soc.spi_video_ram_1.write_fifo.fifo_mem\[30\]\[12\] _04011_ _04014_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_243_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_188_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09598_ soc.rom_encoder_0.input_buffer\[7\] _04600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_184_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08549_ _02138_ soc.spi_video_ram_1.write_fifo.fifo_mem\[2\]\[9\] _03967_ _03977_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_93_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_126_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_208_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11560_ _00626_ clknet_leaf_231_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[25\]\[25\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_243_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_196_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10511_ _05015_ _05019_ _05223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_210_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11491_ _00557_ clknet_leaf_318_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[24\]\[14\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_221_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10442_ _05166_ _05167_ _05168_ _02539_ _05169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XFILLER_40_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xcaravel_hack_soc_101 io_oeb[14] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xcaravel_hack_soc_112 io_out[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_137_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xcaravel_hack_soc_123 io_out[32] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_136_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xcaravel_hack_soc_134 la_data_out[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xcaravel_hack_soc_145 la_data_out[17] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_200_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10373_ _02223_ soc.spi_video_ram_1.write_fifo.fifo_mem\[6\]\[3\] _05124_ _05128_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xcaravel_hack_soc_156 la_data_out[29] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_3_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xcaravel_hack_soc_167 la_data_out[40] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xcaravel_hack_soc_178 la_data_out[51] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_152_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12112_ _01140_ clknet_leaf_266_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[6\]\[4\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xcaravel_hack_soc_189 la_data_out[62] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_12043_ net20 clknet_leaf_297_wb_clk_i soc.rom_encoder_0.data_out\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_219_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_151_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_49_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_218_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3140 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3151 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3162 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_46_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3173 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_206_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3184 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_233_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11827_ _00886_ clknet_leaf_102_wb_clk_i soc.rom_encoder_0.input_buffer\[1\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_18_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1760 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1771 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1782 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_230_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1793 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11758_ _00819_ clknet_leaf_61_wb_clk_i soc.spi_video_ram_1.state_sram_clk_counter\[1\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffnq_2
XFILLER_144_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_202_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_1284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10709_ _03563_ _05324_ _05335_ _01267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_179_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11689_ _00750_ clknet_leaf_145_wb_clk_i soc.spi_video_ram_1.fifo_in_data\[7\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_70_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_196_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_216_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07920_ soc.spi_video_ram_1.write_fifo.fifo_mem\[29\]\[21\] _03563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_69_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_155_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_190_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_151_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07851_ _03139_ _03494_ _03495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_25_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_140_wb_clk_i clknet_5_25_0_wb_clk_i clknet_leaf_140_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_06802_ _02477_ soc.ram_encoder_0.output_bits_left\[2\] _02478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_28_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_56_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07782_ _02920_ soc.spi_video_ram_1.write_fifo.fifo_mem\[17\]\[23\] _03427_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xinput2 io_in[11] net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_110_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_237_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09521_ _04545_ _00869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06733_ _02422_ _00204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_209_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_227_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09452_ _04499_ _02525_ _03767_ soc.rom_encoder_0.request_data_out\[8\] _04500_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_149_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_225_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06664_ _02163_ soc.spi_video_ram_1.write_fifo.fifo_mem\[12\]\[21\] _02356_ _02380_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_25_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_08403_ _03897_ _03898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_05615_ soc.spi_video_ram_1.output_buffer\[12\] soc.spi_video_ram_1.output_buffer\[13\]
+ _01468_ _01524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_196_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09383_ _01387_ _04449_ _04450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_40_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06595_ soc.spi_video_ram_1.write_fifo.fifo_mem\[13\]\[19\] _02341_ _02328_ _02342_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_33_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_162_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_33_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08334_ _02175_ soc.spi_video_ram_1.write_fifo.fifo_mem\[1\]\[27\] _03830_ _03860_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_127_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05546_ soc.cpu.AReg.data\[13\] _01456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_71_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_221_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08265_ _02479_ _02493_ _03821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_14_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05477_ _01385_ _01392_ _01393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07216_ _02596_ _02867_ _02618_ _02868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08196_ _02442_ _02463_ _03765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_118_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07147_ soc.spi_video_ram_1.write_fifo.fifo_mem\[8\]\[5\] soc.spi_video_ram_1.write_fifo.fifo_mem\[9\]\[5\]
+ soc.spi_video_ram_1.write_fifo.fifo_mem\[10\]\[5\] soc.spi_video_ram_1.write_fifo.fifo_mem\[11\]\[5\]
+ _02635_ _02636_ _02802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
Xclkbuf_leaf_299_wb_clk_i clknet_5_1_0_wb_clk_i clknet_leaf_299_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_49_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_238_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07078_ _02670_ _02676_ _02733_ _02735_ _00235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
Xclkbuf_leaf_228_wb_clk_i clknet_5_20_0_wb_clk_i clknet_leaf_228_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_117_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06029_ _01916_ _01918_ _01922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_120_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_102_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_101_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09719_ soc.ram_encoder_0.initializing_step\[1\] soc.ram_encoder_0.initializing_step\[0\]
+ _04684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_60_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10991_ _00057_ clknet_leaf_76_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[17\]\[16\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_27_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_16_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_4_6_0_wb_clk_i clknet_3_3_0_wb_clk_i clknet_4_6_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_245_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_43_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_215_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_150_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11612_ _00678_ clknet_leaf_31_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[21\]\[19\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_212_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_180_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11543_ _00609_ clknet_5_29_0_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[25\]\[8\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_129_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_211_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11474_ _00540_ clknet_leaf_281_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[15\]\[26\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_184_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_193_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10425_ _05154_ _01164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_67_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_100_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_217_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_193_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10356_ soc.cpu.ALU.x\[12\] _05109_ _05118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_98_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_140_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_174_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10287_ soc.rom_loader.current_address\[1\] _05069_ soc.rom_loader.current_address\[2\]
+ _05075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_183_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_1474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12026_ _01085_ clknet_leaf_313_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[5\]\[14\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_191_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_1428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_238_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_219_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_207_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_185_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_146_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_221_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_1286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_33_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_146_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06380_ _02208_ _00065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_203_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_179_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_147_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08050_ soc.spi_video_ram_1.write_fifo.fifo_mem\[11\]\[3\] _02397_ _03680_ _03684_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_204_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07001_ _02583_ _02660_ _02640_ _02661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_190_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_116_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_239_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_321_wb_clk_i clknet_5_0_0_wb_clk_i clknet_leaf_321_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_102_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08952_ _04197_ _00647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_115_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07903_ _02952_ _03543_ _03545_ _03546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_08883_ _04160_ _00615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_29_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07834_ _03047_ soc.spi_video_ram_1.write_fifo.fifo_mem\[17\]\[22\] _03478_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_170_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3909 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07765_ soc.spi_video_ram_1.write_fifo.fifo_mem\[9\]\[15\] _03410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_84_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06716_ _02413_ _00196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09504_ _02258_ soc.cpu.AReg.data\[4\] _04339_ _04537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_246_1626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07696_ _02601_ _03341_ _03342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_52_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_164_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09435_ soc.rom_encoder_0.request_data_out\[4\] _03767_ _04487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_73_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06647_ _02371_ _00169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_197_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_94_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_36_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09366_ _04437_ _04438_ _00820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_36_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06578_ _02331_ _00140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_244_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_240_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_184_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_166_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08317_ _03851_ _00358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05529_ soc.spi_video_ram_1.initialized _00010_ _01440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_166_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09297_ _02223_ soc.spi_video_ram_1.write_fifo.fifo_mem\[4\]\[3\] _04395_ _04399_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_201_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_222_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08248_ _02558_ _03806_ _03807_ _00333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_123_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_197_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_opt_1_0_wb_clk_i clknet_5_10_0_wb_clk_i clknet_opt_1_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_21_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08179_ _03755_ _00316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_175_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10210_ _02219_ soc.spi_video_ram_1.write_fifo.fifo_mem\[5\]\[1\] _05030_ _05032_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_88_1474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_137_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11190_ _00256_ clknet_leaf_191_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[11\]\[0\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_6502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10141_ soc.ram_data_out\[14\] _04928_ _04981_ _04982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_134_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5801 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5812 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_88_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5823 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10072_ _04926_ _04927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_6579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5834 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_173_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5845 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_198_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5856 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_5867 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5878 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5889 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_210_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10974_ _00040_ clknet_leaf_303_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[18\]\[28\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_44_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_244_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_203_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_147_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_176_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_169_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_180_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11526_ _00592_ clknet_leaf_50_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[23\]\[20\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_102_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11457_ _00523_ clknet_leaf_257_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[15\]\[9\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10408_ _02258_ soc.spi_video_ram_1.write_fifo.fifo_mem\[6\]\[20\] _05123_ _05146_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_11388_ _00454_ clknet_leaf_272_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[28\]\[27\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_139_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10339_ _05102_ _05109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_140_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_61_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_234_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12009_ _01068_ clknet_leaf_163_wb_clk_i soc.hack_clock_0.counter\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_05880_ _01669_ _01776_ _01777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_66_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_187_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07550_ _02693_ _03193_ _03196_ _02984_ _03197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_228_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06501_ _02136_ soc.spi_video_ram_1.write_fifo.fifo_mem\[0\]\[8\] _02279_ _02288_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_165_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_234_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_179_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07481_ _02919_ _03128_ _03129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09220_ _04052_ _04346_ _04356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_50_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06432_ _02243_ _00082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_195_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_222_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09151_ soc.spi_video_ram_1.state_counter\[10\] _04311_ _04312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_06363_ _02153_ soc.spi_video_ram_1.write_fifo.fifo_mem\[17\]\[16\] _02193_ _02200_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_175_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08102_ _03710_ _00284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_175_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09082_ _04271_ _00703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06294_ _02157_ soc.spi_video_ram_1.write_fifo.fifo_mem\[18\]\[18\] _02141_ _02158_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_148_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_194_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08033_ _02768_ _03670_ _03671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_162_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_1753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_103_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09984_ _02484_ _02486_ _04873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_103_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5108 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5119 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08935_ _04188_ _00639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_69_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08866_ _04151_ _00607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_131_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3706 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_244_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3717 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_57_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07817_ _02752_ soc.spi_video_ram_1.write_fifo.fifo_mem\[8\]\[23\] _03461_ _03462_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_3728 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3739 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08797_ _04114_ _00575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07748_ soc.spi_video_ram_1.write_fifo.fifo_mem\[31\]\[15\] _03393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_26_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_232_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_226_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_246_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_77_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07679_ _02574_ soc.spi_video_ram_1.write_fifo.fifo_mem\[6\]\[14\] _03324_ _02894_
+ _03325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_38_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_201_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09418_ soc.rom_encoder_0.request_data_out\[0\] _03767_ _04474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_10690_ soc.spi_video_ram_1.fifo_in_data\[12\] _05325_ _05326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_40_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_1530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_205_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_185_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_179_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09349_ _04425_ _00816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_142_1443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_194_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_243_wb_clk_i clknet_5_17_0_wb_clk_i clknet_leaf_243_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_240_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11311_ _00377_ clknet_leaf_184_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[26\]\[8\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_14_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_181_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12291_ _01319_ clknet_leaf_312_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[7\]\[15\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_14_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11242_ _00308_ clknet_leaf_12_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[10\]\[13\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_84_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_84_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_218_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_136_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11173_ _00239_ clknet_leaf_56_wb_clk_i soc.spi_video_ram_1.output_buffer\[17\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_6321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_231_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10124_ _04861_ _04947_ _04948_ _04968_ _04969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_6354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_118_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_212_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_236_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10055_ _04913_ _01035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_231_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4930 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4941 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_5686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5697 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4952 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4963 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4974 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4985 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_169_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4996 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_169_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_229_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_189_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_216_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xclkbuf_5_15_0_wb_clk_i clknet_4_7_0_wb_clk_i clknet_5_15_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_10957_ _00023_ clknet_leaf_33_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[18\]\[11\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_90_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_204_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10888_ _05432_ _01349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_148_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_160_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_8_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_195_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11509_ _00575_ clknet_leaf_134_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[23\]\[3\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12489_ net49 net47 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_176_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_160_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_140_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06981_ _02571_ _02639_ _02640_ _02641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_224_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_86_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05932_ _01822_ _01825_ _01826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_6_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08720_ soc.spi_video_ram_1.write_fifo.fifo_mem\[15\]\[27\] _02351_ _04043_ _04072_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xclkbuf_leaf_47_wb_clk_i clknet_5_9_0_wb_clk_i clknet_leaf_47_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_117_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_226_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08651_ _04030_ _00513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_39_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05863_ _01561_ _01760_ _01761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_94_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_242_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07602_ soc.spi_video_ram_1.write_fifo.fifo_mem\[29\]\[25\] _03249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_54_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08582_ _02171_ soc.spi_video_ram_1.write_fifo.fifo_mem\[2\]\[25\] _03966_ _03994_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_214_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_208_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05794_ _01684_ _01688_ _01696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07533_ _02706_ _03177_ _03180_ _03181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_74_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_241_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_208_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07464_ soc.spi_video_ram_1.write_fifo.fifo_mem\[21\]\[12\] _03112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_224_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09203_ _00011_ _01680_ _04347_ _00748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06415_ soc.spi_video_ram_1.write_fifo.fifo_mem\[16\]\[7\] _02231_ _02217_ _02232_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_72_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07395_ _02926_ soc.spi_video_ram_1.write_fifo.fifo_mem\[12\]\[11\] _03044_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_202_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_194_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09134_ soc.spi_video_ram_1.state_counter\[4\] _04298_ _04301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_148_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06346_ _02136_ soc.spi_video_ram_1.write_fifo.fifo_mem\[17\]\[8\] _02182_ _02191_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_147_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_198_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09065_ _04262_ _00695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_163_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06277_ _02146_ _00024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_191_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08016_ _03645_ _03654_ _03655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_85_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_235_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09967_ soc.ram_encoder_0.input_buffer\[2\] _04849_ _04248_ _04862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_134_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_213_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_131_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_4204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_218_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08918_ soc.spi_video_ram_1.write_fifo.fifo_mem\[22\]\[1\] _02393_ _04178_ _04180_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_09898_ _02454_ _04810_ _04601_ _04811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_4226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08849_ _04141_ _00600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_100_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2802 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_84_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2813 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11860_ _00919_ clknet_leaf_106_wb_clk_i soc.rom_encoder_0.request_address\[5\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2824 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_233_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2835 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2846 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2857 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10811_ _05390_ _01314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_11791_ _00852_ clknet_leaf_130_wb_clk_i soc.spi_video_ram_1.buffer_index\[2\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_2_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2868 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_198_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2879 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10742_ soc.spi_video_ram_1.write_fifo.fifo_mem\[31\]\[8\] soc.spi_video_ram_1.fifo_in_data\[8\]
+ _05344_ _05353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_246_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_230_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10673_ _02227_ soc.spi_video_ram_1.write_fifo.fifo_mem\[29\]\[5\] _05310_ _05316_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_142_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_1314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12343_ _01371_ clknet_leaf_252_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[8\]\[22\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_86_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_182_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_142_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12274_ _01302_ clknet_leaf_270_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[31\]\[27\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_5_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11225_ _00291_ clknet_leaf_87_wb_clk_i soc.video_generator_1.h_count\[6\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_4_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_190_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11156_ _00222_ clknet_leaf_93_wb_clk_i soc.rom_encoder_0.output_bits_left\[3\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_150_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6140 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6151 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6162 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_7_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6173 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10107_ soc.ram_encoder_0.request_data_out\[6\] _04930_ _04956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6184 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_136_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_5450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_191_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11087_ _00153_ clknet_leaf_285_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[13\]\[25\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_237_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_49_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_208_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10038_ soc.ram_encoder_0.request_address\[5\] soc.ram_encoder_0.address\[5\] _04900_
+ _04905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_97_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4760 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4771 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_224_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_188_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4782 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4793 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_223_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_16_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11989_ _01048_ clknet_leaf_118_wb_clk_i soc.ram_data_out\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_182_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_220_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_225_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_165_wb_clk_i clknet_5_30_0_wb_clk_i clknet_leaf_165_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_127_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_182_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06200_ _02086_ net71 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_176_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_203_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_160_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07180_ soc.spi_video_ram_1.write_fifo.fifo_mem\[0\]\[6\] soc.spi_video_ram_1.write_fifo.fifo_mem\[1\]\[6\]
+ soc.spi_video_ram_1.write_fifo.fifo_mem\[2\]\[6\] soc.spi_video_ram_1.write_fifo.fifo_mem\[3\]\[6\]
+ _02613_ _02652_ _02834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_76_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_129_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_199_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06131_ _01955_ _01956_ _02024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_8_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06062_ _01848_ _01890_ _01955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_126_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_232_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_235_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09821_ soc.cpu.DMuxJMP.sel\[1\] _04740_ _04750_ _04751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_28_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09752_ _04705_ _00940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06964_ _01419_ _02624_ _02625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_80_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_100_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_227_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08703_ soc.spi_video_ram_1.fifo_in_address\[5\] _04061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_05915_ _01705_ _01809_ _01810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_104_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09683_ soc.cpu.PC.REG.data\[7\] _04656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_06895_ _02556_ _02557_ _02559_ _00229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_94_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2109 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_243_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05846_ _01740_ _01743_ _01745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_08634_ _02161_ soc.spi_video_ram_1.write_fifo.fifo_mem\[30\]\[20\] _03999_ _04022_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_94_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_215_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05777_ _01615_ _01668_ _01679_ _01680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
X_08565_ _03985_ _00472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_35_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_243_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07516_ _02707_ _03156_ _03163_ _02970_ _03164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_08496_ _02147_ soc.spi_video_ram_1.write_fifo.fifo_mem\[28\]\[13\] _03945_ _03949_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_180_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_1284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_210_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07447_ _02924_ soc.spi_video_ram_1.write_fifo.fifo_mem\[30\]\[27\] _02827_ _03096_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_74_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07378_ _02784_ soc.spi_video_ram_1.write_fifo.fifo_mem\[22\]\[11\] _03027_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_221_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09117_ _02274_ soc.spi_video_ram_1.write_fifo.fifo_mem\[20\]\[28\] _04258_ _04289_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06329_ _02181_ _02182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_108_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_30_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_159_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_104_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_178_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09048_ soc.spi_video_ram_1.write_fifo.read_pointer\[2\] _04247_ _04251_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_124_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_190_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11010_ _00076_ clknet_leaf_211_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[16\]\[6\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_145_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_131_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_219_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4001 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4012 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4023 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4034 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4045 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_180_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4056 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4067 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_206_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4078 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_4089 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11912_ _00971_ clknet_5_13_0_wb_clk_i soc.cpu.ALU.ny vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_205_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11843_ _00902_ clknet_leaf_95_wb_clk_i soc.rom_encoder_0.request_data_out\[4\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1920 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_199_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1942 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_202_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_183_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_246_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1953 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2698 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11774_ _00835_ clknet_leaf_105_wb_clk_i soc.rom_encoder_0.output_buffer\[5\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1964 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1975 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1986 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_207_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_186_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1997 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10725_ _05343_ _05344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_201_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_174_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10656_ _05306_ _01243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_10_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_196_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10587_ _05267_ _05268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_6_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12326_ _01354_ clknet_leaf_189_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[8\]\[5\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_138_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12257_ _01285_ clknet_leaf_13_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[31\]\[10\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_155_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_233_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11208_ _00274_ clknet_leaf_25_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[11\]\[18\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_123_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12188_ _01216_ net87 soc.gpio_i_stored\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_155_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11139_ _00205_ clknet_leaf_28_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[14\]\[19\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_209_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_42_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_49_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05700_ _01598_ soc.cpu.AReg.data\[1\] _01600_ _01605_ _01606_ _01607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
XFILLER_3_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_225_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_149_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06680_ soc.spi_video_ram_1.write_fifo.write_pointer\[1\] _01444_ _02388_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_4590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_52_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05631_ _01468_ soc.spi_video_ram_1.output_buffer\[5\] _01540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_36_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08350_ _03870_ _00372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05562_ _01469_ _01470_ _01471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_189_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_244_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07301_ _02949_ _02950_ _02598_ _02951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_08281_ _02122_ soc.spi_video_ram_1.write_fifo.fifo_mem\[1\]\[1\] _03831_ _03833_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_162_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05493_ _01402_ _01404_ _01406_ _01407_ _01408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_53_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_123_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07232_ _02883_ _00241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_165_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_101_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_9_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07163_ _02650_ _02817_ _02618_ _02818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_9_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06114_ _01967_ _01988_ _01986_ _02007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_117_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_238_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_172_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07094_ _02726_ soc.spi_video_ram_1.write_fifo.fifo_mem\[14\]\[3\] _02714_ _02751_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xclkbuf_5_8_0_wb_clk_i clknet_4_4_0_wb_clk_i clknet_5_8_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_195_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06045_ _01896_ _01936_ _01937_ _01934_ _01938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
Xclkbuf_leaf_62_wb_clk_i clknet_5_12_0_wb_clk_i clknet_leaf_62_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_236_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09804_ _01396_ _04735_ _00962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_41_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07996_ soc.spi_video_ram_1.output_buffer\[3\] _02676_ _03636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_45_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_1745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09735_ _04695_ _04696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_41_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06947_ soc.spi_video_ram_1.write_fifo.fifo_mem\[28\]\[0\] soc.spi_video_ram_1.write_fifo.fifo_mem\[29\]\[0\]
+ soc.spi_video_ram_1.write_fifo.fifo_mem\[30\]\[0\] soc.spi_video_ram_1.write_fifo.fifo_mem\[31\]\[0\]
+ _02607_ _02578_ _02608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_55_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09666_ soc.cpu.PC.REG.data\[2\] soc.rom_loader.current_address\[2\] _04638_ _04644_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06878_ _02545_ _00226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_41_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08617_ _04013_ _00496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_83_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_242_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05829_ _01716_ _01721_ _01729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09597_ _04598_ _04585_ _04599_ _00891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_110_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08548_ _03976_ _00464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_51_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_211_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08479_ _02130_ soc.spi_video_ram_1.write_fifo.fifo_mem\[28\]\[5\] _03934_ _03940_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_145_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10510_ _05221_ _05222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_50_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_11490_ _00556_ clknet_leaf_314_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[24\]\[13\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_126_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10441_ _01779_ _01819_ _05163_ _05168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
Xcaravel_hack_soc_102 io_oeb[15] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xcaravel_hack_soc_113 io_out[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xcaravel_hack_soc_124 io_out[33] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xcaravel_hack_soc_135 la_data_out[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_137_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10372_ _05127_ _01138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xcaravel_hack_soc_146 la_data_out[18] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_139_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_191_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xcaravel_hack_soc_157 la_data_out[30] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xcaravel_hack_soc_168 la_data_out[41] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_163_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12111_ _01139_ clknet_leaf_266_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[6\]\[3\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xcaravel_hack_soc_179 la_data_out[52] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_46_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12042_ _01101_ clknet_leaf_125_wb_clk_i soc.rom_loader.writing vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_46_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_238_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_213_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_207_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3130 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3141 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3152 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_234_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3163 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3174 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3185 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11826_ _00885_ clknet_leaf_125_wb_clk_i soc.rom_encoder_0.input_buffer\[0\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1750 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1761 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_226_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1772 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1783 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1794 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11757_ _00818_ clknet_leaf_61_wb_clk_i soc.spi_video_ram_1.state_sram_clk_counter\[0\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffnq_2
XFILLER_197_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_159_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_204_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_140_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10708_ soc.spi_video_ram_1.fifo_in_address\[5\] _05325_ _05335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_105_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11688_ _00749_ clknet_leaf_145_wb_clk_i soc.spi_video_ram_1.fifo_in_data\[6\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_220_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_161_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10639_ soc.spi_video_ram_1.write_fifo.fifo_mem\[19\]\[18\] soc.spi_video_ram_1.fifo_in_address\[2\]
+ _05289_ _05298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_143_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12309_ _01337_ clknet_leaf_155_wb_clk_i soc.ram_encoder_0.data_out\[4\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_237_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07850_ soc.spi_video_ram_1.write_fifo.fifo_mem\[29\]\[22\] _03494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_96_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06801_ soc.ram_encoder_0.output_bits_left\[3\] _02477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_7_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_232_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07781_ soc.spi_video_ram_1.write_fifo.fifo_mem\[18\]\[23\] soc.spi_video_ram_1.write_fifo.fifo_mem\[19\]\[23\]
+ _02591_ _03426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_83_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xinput3 io_in[12] net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_37_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09520_ _02274_ soc.cpu.AReg.data\[12\] _01459_ _04545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06732_ soc.spi_video_ram_1.write_fifo.fifo_mem\[14\]\[18\] _02339_ _02412_ _02422_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_37_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_180_wb_clk_i clknet_5_29_0_wb_clk_i clknet_leaf_180_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_52_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09451_ soc.rom_encoder_0.request_write _04499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_65_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06663_ _02379_ _00177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_224_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08402_ _01441_ _03863_ _03897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05614_ _01469_ _01518_ _01523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_244_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06594_ soc.spi_video_ram_1.fifo_in_address\[3\] _02341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_09382_ soc.spi_video_ram_1.state_sram_clk_counter\[7\] _04445_ _04449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_240_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_178_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05545_ soc.cpu.instruction\[15\] soc.cpu.instruction\[3\] _01455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_08333_ _03859_ _00366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_71_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_220_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08264_ _03820_ _00336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_32_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05476_ _01386_ _01391_ _01392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_07215_ soc.spi_video_ram_1.write_fifo.fifo_mem\[4\]\[8\] soc.spi_video_ram_1.write_fifo.fifo_mem\[5\]\[8\]
+ soc.spi_video_ram_1.write_fifo.fifo_mem\[6\]\[8\] soc.spi_video_ram_1.write_fifo.fifo_mem\[7\]\[8\]
+ _02597_ _02598_ _02867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_193_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08195_ _03763_ _02458_ _03764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_203_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07146_ _01508_ _02676_ _02735_ _02801_ _00237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_140_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_192_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_3_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07077_ _01409_ _01411_ _02734_ _02626_ _02735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_82_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06028_ _01848_ _01890_ _01920_ _01921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_82_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_216_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_268_wb_clk_i clknet_5_7_0_wb_clk_i clknet_leaf_268_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_134_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_60_1520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07979_ soc.spi_video_ram_1.write_fifo.fifo_mem\[12\]\[18\] soc.spi_video_ram_1.write_fifo.fifo_mem\[13\]\[18\]
+ soc.spi_video_ram_1.write_fifo.fifo_mem\[14\]\[18\] soc.spi_video_ram_1.write_fifo.fifo_mem\[15\]\[18\]
+ _02726_ _03041_ _03619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_169_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_210_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09718_ soc.ram_encoder_0.initializing_step\[2\] _04683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_10990_ _00056_ clknet_leaf_10_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[17\]\[15\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_216_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09649_ _04633_ _00909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_243_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_1728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_180_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11611_ _00677_ clknet_leaf_28_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[21\]\[18\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_208_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_169_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_243_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_196_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11542_ _00608_ clknet_leaf_146_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[25\]\[7\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_11_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_221_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11473_ _00539_ clknet_leaf_285_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[15\]\[25\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_87_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10424_ _02274_ soc.spi_video_ram_1.write_fifo.fifo_mem\[6\]\[28\] _05123_ _05154_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_139_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10355_ _01779_ _05104_ _05117_ _01131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_124_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_234_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10286_ _05074_ _01104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_219_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_152_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_156_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12025_ _01084_ clknet_leaf_312_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[5\]\[13\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_239_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_65_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_202_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_206_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_185_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_222_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_146_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11809_ _00869_ clknet_leaf_270_wb_clk_i soc.spi_video_ram_1.fifo_in_address\[12\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_241_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_221_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_202_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_1468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_187_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_109_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_186_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_70_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07000_ soc.spi_video_ram_1.write_fifo.fifo_mem\[24\]\[1\] soc.spi_video_ram_1.write_fifo.fifo_mem\[25\]\[1\]
+ soc.spi_video_ram_1.write_fifo.fifo_mem\[26\]\[1\] soc.spi_video_ram_1.write_fifo.fifo_mem\[27\]\[1\]
+ _02635_ _02636_ _02660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_122_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_200_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_179_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_157_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_227_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_196_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08951_ soc.spi_video_ram_1.write_fifo.fifo_mem\[22\]\[17\] _02337_ _04189_ _04197_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_174_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07902_ _02704_ soc.spi_video_ram_1.write_fifo.fifo_mem\[13\]\[21\] _03544_ _02742_
+ _03545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_29_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08882_ soc.spi_video_ram_1.write_fifo.fifo_mem\[25\]\[14\] _04052_ _04155_ _04160_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_57_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_233_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_243_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_229_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07833_ soc.spi_video_ram_1.write_fifo.fifo_mem\[18\]\[22\] soc.spi_video_ram_1.write_fifo.fifo_mem\[19\]\[22\]
+ _02575_ _03477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_42_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_211_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07764_ _02922_ soc.spi_video_ram_1.write_fifo.fifo_mem\[11\]\[15\] _02647_ _03409_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09503_ _04536_ _00860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06715_ soc.spi_video_ram_1.write_fifo.fifo_mem\[14\]\[10\] _02411_ _02412_ _02413_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_112_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_225_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07695_ _02900_ _03337_ _03340_ _03341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_24_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09434_ _04473_ _04485_ _04486_ _00841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_20_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06646_ _02145_ soc.spi_video_ram_1.write_fifo.fifo_mem\[12\]\[12\] _02368_ _02371_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XPHY_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_164_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_1697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09365_ soc.spi_video_ram_1.state_sram_clk_counter\[2\] _04435_ _04433_ _04438_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06577_ soc.spi_video_ram_1.write_fifo.fifo_mem\[13\]\[12\] _02242_ _02328_ _02331_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_209_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_221_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08316_ _02157_ soc.spi_video_ram_1.write_fifo.fifo_mem\[1\]\[18\] _03842_ _03851_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_240_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05528_ _01439_ _00010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_55_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09296_ _04398_ _00790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08247_ soc.ram_encoder_0.output_buffer\[13\] _02555_ _03807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_181_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08178_ _02163_ soc.spi_video_ram_1.write_fifo.fifo_mem\[10\]\[21\] _03731_ _03755_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_146_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07129_ _02784_ soc.spi_video_ram_1.write_fifo.fifo_mem\[13\]\[4\] _02785_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_238_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_84_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10140_ _04869_ _04930_ _04926_ _04980_ _04981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_6514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_133_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5802 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5813 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10071_ _02480_ _02481_ _04925_ _04926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XTAP_6569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5824 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5835 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5846 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5857 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_102_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5868 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_47_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_1749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5879 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_169_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_16_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10973_ _00039_ clknet_leaf_271_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[18\]\[27\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_189_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_43_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_204_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_186_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_203_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_197_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_200_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11525_ _00591_ clknet_leaf_32_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[23\]\[19\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_89_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_141_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_184_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_172_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11456_ _00522_ clknet_leaf_177_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[15\]\[8\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_67_1515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10407_ _05145_ _01155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_217_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11387_ _00453_ clknet_leaf_294_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[28\]\[26\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_98_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_180_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10338_ _01652_ _05103_ _05108_ _01123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_119_wb_clk_i clknet_5_26_0_wb_clk_i clknet_leaf_119_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_139_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_191_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10269_ soc.rom_encoder_0.initialized _04611_ _05063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_117_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12008_ _01067_ clknet_leaf_163_wb_clk_i soc.hack_clock_0.counter\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_121_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_238_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_207_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06500_ _02287_ _00106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07480_ soc.spi_video_ram_1.write_fifo.fifo_mem\[5\]\[12\] _03128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_146_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_228_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06431_ soc.spi_video_ram_1.write_fifo.fifo_mem\[16\]\[12\] _02242_ _02238_ _02243_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_188_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_203_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09150_ soc.spi_video_ram_1.state_counter\[9\] _04308_ _04311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06362_ _02199_ _00056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_175_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_241_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_187_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08101_ soc.spi_video_ram_1.write_fifo.fifo_mem\[11\]\[28\] _02353_ _03679_ _03710_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_09081_ _02237_ soc.spi_video_ram_1.write_fifo.fifo_mem\[20\]\[10\] _04270_ _04271_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06293_ soc.spi_video_ram_1.fifo_in_address\[2\] _02157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_190_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08032_ soc.spi_video_ram_1.write_fifo.fifo_mem\[16\]\[16\] soc.spi_video_ram_1.write_fifo.fifo_mem\[17\]\[16\]
+ soc.spi_video_ram_1.write_fifo.fifo_mem\[18\]\[16\] soc.spi_video_ram_1.write_fifo.fifo_mem\[19\]\[16\]
+ _02681_ _02758_ _03670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_116_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_239_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09983_ _04871_ _04849_ _04872_ _01004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_89_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_170_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5109 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08934_ soc.spi_video_ram_1.write_fifo.fifo_mem\[22\]\[9\] _02409_ _04178_ _04188_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_192_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_1353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_4408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08865_ soc.spi_video_ram_1.write_fifo.fifo_mem\[25\]\[6\] _02403_ _04144_ _04151_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_170_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3707 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07816_ _02763_ _03460_ _03461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_3718 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3729 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08796_ _02126_ soc.spi_video_ram_1.write_fifo.fifo_mem\[23\]\[3\] _04110_ _04114_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_246_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07747_ soc.spi_video_ram_1.write_fifo.fifo_mem\[24\]\[15\] soc.spi_video_ram_1.write_fifo.fifo_mem\[25\]\[15\]
+ soc.spi_video_ram_1.write_fifo.fifo_mem\[26\]\[15\] soc.spi_video_ram_1.write_fifo.fifo_mem\[27\]\[15\]
+ _02688_ _02827_ _03392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_244_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_183_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_16_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_164_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07678_ _02902_ _03323_ _03324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_207_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_197_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09417_ _02541_ _04473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_13_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06629_ _02128_ soc.spi_video_ram_1.write_fifo.fifo_mem\[12\]\[4\] _02357_ _02362_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_129_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_244_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_240_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_199_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09348_ _02274_ soc.spi_video_ram_1.write_fifo.fifo_mem\[4\]\[28\] _04394_ _04425_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_181_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09279_ _04069_ _04360_ _04388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_166_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11310_ _00376_ clknet_leaf_146_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[26\]\[7\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_138_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12290_ _01318_ clknet_leaf_312_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[7\]\[14\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_119_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11241_ _00307_ clknet_leaf_1_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[10\]\[12\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_106_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_175_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_1242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_283_wb_clk_i clknet_5_7_0_wb_clk_i clknet_leaf_283_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_10_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_162_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11172_ _00238_ clknet_leaf_55_wb_clk_i soc.spi_video_ram_1.output_buffer\[18\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_6311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_175_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_175_1286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_212_wb_clk_i clknet_5_20_0_wb_clk_i clknet_leaf_212_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_6333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10123_ soc.ram_encoder_0.request_data_out\[10\] _04929_ _04968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_6344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10054_ soc.ram_encoder_0.request_address\[13\] soc.ram_encoder_0.address\[13\] _04879_
+ _04913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_5654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_6399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4920 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4931 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4942 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5698 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4953 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4964 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_236_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4975 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4986 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4997 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_56_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10956_ _00022_ clknet_leaf_18_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[18\]\[10\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_147_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_229_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_232_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10887_ soc.spi_video_ram_1.write_fifo.fifo_mem\[8\]\[0\] soc.spi_video_ram_1.fifo_in_data\[0\]
+ _05431_ _05432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XPHY_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_34_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_199_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11508_ _00574_ clknet_leaf_55_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[23\]\[2\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12488_ net49 net46 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_145_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11439_ _00505_ clknet_leaf_49_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[30\]\[20\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_158_1451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_1501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06980_ _02585_ _02640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_26_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_234_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05931_ _01705_ _01824_ _01825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_26_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_113_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_239_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08650_ _02177_ soc.spi_video_ram_1.write_fifo.fifo_mem\[30\]\[28\] _03999_ _04030_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_05862_ _01717_ _01759_ _01760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_212_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_187_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07601_ _02575_ soc.spi_video_ram_1.write_fifo.fifo_mem\[30\]\[25\] _03247_ _02904_
+ _03248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_08581_ _03993_ _00480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_240_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_87_wb_clk_i clknet_5_11_0_wb_clk_i clknet_leaf_87_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_05793_ _01689_ _01694_ _01695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_226_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07532_ _02700_ soc.spi_video_ram_1.write_fifo.fifo_mem\[4\]\[26\] _03179_ _02741_
+ _03180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_81_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_165_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_179_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_16_wb_clk_i clknet_5_2_0_wb_clk_i clknet_leaf_16_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_23_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07463_ _02607_ soc.spi_video_ram_1.write_fifo.fifo_mem\[22\]\[12\] _03110_ _02904_
+ _03111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_195_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_222_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09202_ soc.spi_video_ram_1.fifo_in_data\[5\] _04346_ _04347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_245_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06414_ soc.spi_video_ram_1.fifo_in_data\[7\] _02231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_07394_ _02920_ soc.spi_video_ram_1.write_fifo.fifo_mem\[13\]\[11\] _03043_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09133_ soc.spi_video_ram_1.state_counter\[4\] _04298_ _04300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_06345_ _02190_ _00048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_148_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_191_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06276_ _02145_ soc.spi_video_ram_1.write_fifo.fifo_mem\[18\]\[12\] _02141_ _02146_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_09064_ _02221_ soc.spi_video_ram_1.write_fifo.fifo_mem\[20\]\[2\] _04259_ _04262_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_108_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08015_ _03647_ _03649_ _03651_ _03653_ _02568_ _03654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_200_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_150_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_103_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_137_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09966_ soc.ram_encoder_0.input_buffer\[6\] _04861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_77_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08917_ _04179_ _00630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_170_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_4205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09897_ _04573_ _04809_ _04810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_4216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_4227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08848_ _02177_ soc.spi_video_ram_1.write_fifo.fifo_mem\[23\]\[28\] _04109_ _04141_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_57_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_218_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2803 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2814 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08779_ _04103_ _00568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2825 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_232_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_245_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2836 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10810_ _02237_ soc.spi_video_ram_1.write_fifo.fifo_mem\[7\]\[10\] _05389_ _05390_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_2847 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2858 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2869 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11790_ _00851_ clknet_leaf_63_wb_clk_i soc.spi_video_ram_1.buffer_index\[1\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_246_1243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10741_ _05352_ _01282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_214_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_186_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_198_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_185_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10672_ _05315_ _01250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_9_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_1282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_224_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_223_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_154_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12342_ _01370_ clknet_leaf_283_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[8\]\[21\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_127_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_181_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12273_ _01301_ clknet_leaf_294_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[31\]\[26\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_218_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11224_ _00290_ clknet_leaf_86_wb_clk_i soc.video_generator_1.h_count\[5\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_175_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_150_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6130 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11155_ _00221_ clknet_leaf_95_wb_clk_i soc.rom_encoder_0.output_bits_left\[4\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_150_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6141 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_68_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_6152 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_6163 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10106_ _04952_ _04955_ _01043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_6174 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6185 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11086_ _00152_ clknet_leaf_305_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[13\]\[24\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_6196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10037_ _04904_ _01026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_5484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4750 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_114_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_4761 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_237_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4772 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4783 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_208_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4794 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11988_ _01047_ clknet_leaf_158_wb_clk_i soc.ram_data_out\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_147_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_210_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10939_ _05458_ _01374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_32_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_204_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_242_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_220_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06130_ _01921_ _02011_ _02022_ _02023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_144_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_134_wb_clk_i clknet_5_24_0_wb_clk_i clknet_leaf_134_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_145_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06061_ _01927_ _01938_ _01952_ _01954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_173_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_67_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09820_ _04741_ _04748_ _04749_ _04750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_28_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09751_ _02231_ soc.spi_video_ram_1.write_fifo.fifo_mem\[3\]\[7\] _04697_ _04705_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_113_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06963_ soc.spi_video_ram_1.state_sram_clk_counter\[1\] _01391_ _02624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_2
XFILLER_67_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08702_ _04060_ _00534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05914_ _01717_ _01808_ _01809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_132_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09682_ _04468_ _04618_ _04655_ _00920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_39_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06894_ soc.ram_encoder_0.output_buffer\[4\] _02558_ _02559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_82_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08633_ _04021_ _00504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_230_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05845_ _01740_ _01743_ _01744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_110_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_214_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_227_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08564_ _02153_ soc.spi_video_ram_1.write_fifo.fifo_mem\[2\]\[16\] _03978_ _03985_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_05776_ _01669_ _01677_ _01678_ _01679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_74_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_208_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07515_ _02588_ _03159_ _03162_ _03163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_120_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_93_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08495_ _03948_ _00439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_74_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07446_ _02696_ soc.spi_video_ram_1.write_fifo.fifo_mem\[31\]\[27\] _03095_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_161_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_221_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_202_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07377_ _03020_ _03022_ _03023_ _03025_ _02929_ _03026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_136_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09116_ _04288_ _00720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06328_ _02180_ _02181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_163_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_237_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09047_ soc.spi_video_ram_1.write_fifo.read_pointer\[2\] _04247_ _04250_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06259_ soc.spi_video_ram_1.fifo_in_data\[7\] _02134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_159_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_219_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_132_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_77_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_237_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09949_ net1 _04849_ _04601_ _04850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_150_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4002 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4013 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4024 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4035 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4046 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4057 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_219_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4068 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11911_ _00970_ clknet_leaf_127_wb_clk_i soc.cpu.ALU.f vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_4079 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_173_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_233_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11842_ _00901_ clknet_leaf_170_wb_clk_i soc.rom_encoder_0.request_data_out\[3\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_79_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1910 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1921 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1932 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1943 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_220_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11773_ _00834_ clknet_leaf_89_wb_clk_i soc.spi_video_ram_1.read_value\[3\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1954 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2699 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1965 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1976 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1987 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10724_ _01445_ _03931_ _05343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_1998 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_202_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10655_ soc.spi_video_ram_1.write_fifo.fifo_mem\[19\]\[26\] _03927_ _05277_ _05306_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_155_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10586_ _01455_ _01575_ _05267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_155_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_196_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12325_ _01353_ clknet_leaf_197_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[8\]\[4\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_86_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12256_ _01284_ clknet_leaf_257_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[31\]\[9\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_108_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_237_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_64_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_190_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_2_1_0_wb_clk_i clknet_0_wb_clk_i clknet_2_1_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_11207_ _00273_ clknet_leaf_24_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[11\]\[17\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12187_ _01215_ net86 soc.gpio_i_stored\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_229_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_214_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11138_ _00204_ clknet_leaf_22_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[14\]\[18\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_96_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_23_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11069_ _00135_ clknet_leaf_191_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[13\]\[7\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_114_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_95_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_209_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05630_ soc.spi_video_ram_1.output_buffer\[4\] _01539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_3890 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05561_ soc.spi_video_ram_1.buffer_index\[2\] _01470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_75_1466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_225_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07300_ _02941_ soc.spi_video_ram_1.write_fifo.fifo_mem\[16\]\[10\] _02950_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_149_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08280_ _03832_ _00340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05492_ soc.spi_video_ram_1.write_fifo.read_pointer\[4\] soc.spi_video_ram_1.write_fifo.write_pointer\[4\]
+ _01407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
Xclkbuf_leaf_315_wb_clk_i clknet_5_0_0_wb_clk_i clknet_leaf_315_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_07231_ soc.spi_video_ram_1.output_buffer\[15\] _02881_ _02882_ _02883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_203_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_158_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_192_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07162_ soc.spi_video_ram_1.write_fifo.fifo_mem\[20\]\[5\] soc.spi_video_ram_1.write_fifo.fifo_mem\[21\]\[5\]
+ soc.spi_video_ram_1.write_fifo.fifo_mem\[22\]\[5\] soc.spi_video_ram_1.write_fifo.fifo_mem\[23\]\[5\]
+ _02651_ _02652_ _02817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_145_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06113_ _01926_ _02005_ _01967_ _02006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_12_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07093_ _02697_ soc.spi_video_ram_1.write_fifo.fifo_mem\[15\]\[3\] _02750_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_161_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06044_ _01928_ _01929_ _01935_ _01937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_133_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09803_ _04730_ _04734_ soc.rom_encoder_0.initialized _04735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_60_1702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_219_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07995_ _03625_ _03634_ _03635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_74_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09734_ _01445_ _02276_ _04695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06946_ _02590_ _02607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_74_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_31_wb_clk_i clknet_5_9_0_wb_clk_i clknet_leaf_31_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_95_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09665_ _04643_ _00915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_243_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06877_ soc.rom_encoder_0.output_buffer\[3\] _02542_ _02543_ soc.rom_encoder_0.request_address\[2\]
+ _02545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_167_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_215_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08616_ _02143_ soc.spi_video_ram_1.write_fifo.fifo_mem\[30\]\[11\] _04011_ _04013_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_05828_ _01725_ _01727_ _01728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_82_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09596_ soc.rom_encoder_0.input_buffer\[2\] _04586_ _04553_ _04599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_199_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_231_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_243_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_202_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08547_ _02136_ soc.spi_video_ram_1.write_fifo.fifo_mem\[2\]\[8\] _03967_ _03976_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_05759_ _01656_ _01660_ _01663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_196_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08478_ _03939_ _00431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_23_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07429_ _02703_ soc.spi_video_ram_1.write_fifo.fifo_mem\[5\]\[27\] _03078_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_126_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10440_ _01615_ _01833_ _05167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_108_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xcaravel_hack_soc_103 io_oeb[20] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_100_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xcaravel_hack_soc_114 io_out[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xcaravel_hack_soc_125 irq[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_104_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xcaravel_hack_soc_136 la_data_out[8] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_10371_ _02221_ soc.spi_video_ram_1.write_fifo.fifo_mem\[6\]\[2\] _05124_ _05127_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_124_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_164_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xcaravel_hack_soc_147 la_data_out[19] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xcaravel_hack_soc_158 la_data_out[31] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_164_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12110_ _01138_ clknet_leaf_265_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[6\]\[2\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xcaravel_hack_soc_169 la_data_out[42] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_156_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_191_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12041_ _01100_ clknet_leaf_99_wb_clk_i soc.rom_loader.rom_request vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_2_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_215_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3120 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_189_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3131 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3142 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3153 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3164 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3175 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3186 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11825_ _00884_ clknet_leaf_96_wb_clk_i soc.rom_encoder_0.input_bits_left\[4\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_221_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1740 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1751 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1762 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1773 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11756_ _00817_ clknet_leaf_100_wb_clk_i soc.rom_loader.was_loading vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1784 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_222_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_186_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1795 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_201_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10707_ _05334_ _01266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_197_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11687_ _00748_ clknet_leaf_146_wb_clk_i soc.spi_video_ram_1.fifo_in_data\[5\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_128_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10638_ _05297_ _01234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_127_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_196_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10569_ soc.hack_wait_clocks\[0\] _05254_ _05256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_143_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12308_ _01336_ clknet_leaf_155_wb_clk_i soc.ram_encoder_0.data_out\[3\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_5_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12239_ _01267_ clknet_leaf_291_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[29\]\[21\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_233_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06800_ _02453_ _02475_ _02476_ _01381_ _00217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_84_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07780_ _02656_ _03401_ _03424_ _03019_ _03425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_37_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_65_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput4 io_in[13] net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06731_ _02421_ _00203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_225_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09450_ _04473_ _04497_ _04498_ _00845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_64_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06662_ _02161_ soc.spi_video_ram_1.write_fifo.fifo_mem\[12\]\[20\] _02356_ _02379_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_188_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_213_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08401_ _03896_ _00397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05613_ soc.spi_video_ram_1.output_buffer\[14\] soc.spi_video_ram_1.output_buffer\[15\]
+ _01468_ _01522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_09381_ soc.spi_video_ram_1.current_state\[2\] net68 _04448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_06593_ _02340_ _00146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08332_ _02173_ soc.spi_video_ram_1.write_fifo.fifo_mem\[1\]\[26\] _03830_ _03859_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_05544_ soc.hack_wait_clocks\[1\] soc.hack_wait_clocks\[0\] _01452_ _01453_ _01454_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__or4_1
XFILLER_162_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_244_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_177_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08263_ _03819_ soc.ram_encoder_0.output_buffer\[16\] _02555_ _03820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_193_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_20_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05475_ _01387_ soc.spi_video_ram_1.state_sram_clk_counter\[0\] _01390_ _01391_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_119_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07214_ _02589_ _02865_ _02866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_193_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08194_ _02433_ _02437_ _03763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_146_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07145_ _02677_ _02606_ _02791_ _02800_ _02801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_238_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07076_ _02624_ _02671_ _00830_ _02734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_105_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06027_ _01916_ _01918_ _01919_ _01920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_173_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_142_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_28_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07978_ _02736_ _03617_ _03618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09717_ _04680_ _03777_ _03788_ soc.ram_encoder_0.request_data_out\[12\] _04682_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_06929_ _02572_ _02590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_186_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09648_ soc.rom_encoder_0.data_out\[11\] soc.rom_encoder_0.request_data_out\[11\]
+ _04632_ _04633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_95_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_237_wb_clk_i clknet_5_5_0_wb_clk_i clknet_leaf_237_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_110_1390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09579_ _04583_ _04585_ _04587_ _00885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_203_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11610_ _00676_ clknet_leaf_27_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[21\]\[17\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_230_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_168_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_223_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_145_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11541_ _00607_ clknet_leaf_201_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[25\]\[6\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_129_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_156_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11472_ _00538_ clknet_leaf_305_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[15\]\[24\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_109_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_183_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10423_ _05153_ _01163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_109_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_193_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10354_ soc.cpu.ALU.x\[11\] _05109_ _05117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_152_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_174_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10285_ soc.rom_loader.current_address\[1\] _05069_ _05073_ _05074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_140_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12024_ _01083_ clknet_leaf_309_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[5\]\[12\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_234_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_238_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_207_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_234_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_228_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_226_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_241_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_11808_ _00868_ clknet_leaf_263_wb_clk_i soc.spi_video_ram_1.fifo_in_address\[11\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_163_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11739_ _00800_ clknet_leaf_308_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[4\]\[12\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_109_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_239_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_183_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_192_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08950_ _04196_ _00646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_48_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07901_ _02783_ soc.spi_video_ram_1.write_fifo.fifo_mem\[12\]\[21\] _03544_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_97_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08881_ _04159_ _00614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_111_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07832_ _03476_ _00248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_57_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07763_ _02920_ soc.spi_video_ram_1.write_fifo.fifo_mem\[10\]\[15\] _03408_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_186_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09502_ _02256_ soc.cpu.AReg.data\[3\] _04339_ _04536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_71_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06714_ _02389_ _02412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_65_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07694_ _02893_ soc.spi_video_ram_1.write_fifo.fifo_mem\[20\]\[24\] _03339_ _02741_
+ _03340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_65_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_53_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_129_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_246_1639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09433_ soc.rom_encoder_0.output_buffer\[11\] _04479_ _04486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_52_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06645_ _02370_ _00168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_25_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_240_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_212_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09364_ soc.spi_video_ram_1.state_sram_clk_counter\[2\] _04435_ _04437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_24_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06576_ _02330_ _00139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_90_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08315_ _03850_ _00357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05527_ soc.spi_video_ram_1.current_state\[2\] _01412_ _01439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_162_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09295_ _02221_ soc.spi_video_ram_1.write_fifo.fifo_mem\[4\]\[2\] _04395_ _04398_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_123_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08246_ soc.ram_encoder_0.output_buffer\[9\] _03781_ _03789_ soc.ram_encoder_0.request_data_out\[5\]
+ _03805_ _03806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_203_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08177_ _03754_ _00315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_192_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_1443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_10_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07128_ _02783_ _02784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_101_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_6504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_106_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07059_ soc.spi_video_ram_1.write_fifo.fifo_mem\[20\]\[2\] soc.spi_video_ram_1.write_fifo.fifo_mem\[21\]\[2\]
+ soc.spi_video_ram_1.write_fifo.fifo_mem\[22\]\[2\] soc.spi_video_ram_1.write_fifo.fifo_mem\[23\]\[2\]
+ _02717_ _02714_ _02718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_6515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5803 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_216_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10070_ soc.ram_encoder_0.toggled_sram_sck _04924_ _04925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XTAP_6559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5814 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5825 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5836 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5847 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_134_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5858 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_236_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5869 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_130_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_210_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_151_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_216_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_44_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10972_ _00038_ clknet_leaf_288_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[18\]\[26\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_243_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_245_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_227_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_231_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_196_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_169_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11524_ _00590_ clknet_leaf_27_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[23\]\[18\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_12_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11455_ _00521_ clknet_leaf_192_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[15\]\[7\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_165_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10406_ _02256_ soc.spi_video_ram_1.write_fifo.fifo_mem\[6\]\[19\] _05135_ _05145_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_125_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_139_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11386_ _00452_ clknet_leaf_232_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[28\]\[25\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_139_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_193_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10337_ soc.cpu.ALU.x\[3\] _05104_ _05108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_234_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_139_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10268_ _05062_ _01099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_105_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_239_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12007_ _01066_ clknet_leaf_113_wb_clk_i soc.hack_clock_0.counter\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_39_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10199_ soc.hack_clock_0.counter\[4\] _05022_ _05025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_152_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_66_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_159_wb_clk_i clknet_5_27_0_wb_clk_i clknet_leaf_159_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_78_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_235_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_222_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06430_ soc.spi_video_ram_1.fifo_in_data\[12\] _02242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_22_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2090 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06361_ _02151_ soc.spi_video_ram_1.write_fifo.fifo_mem\[17\]\[15\] _02193_ _02199_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_124_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_206_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08100_ _03709_ _00283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_124_1356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09080_ _04257_ _04270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_30_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06292_ _02156_ _00029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_238_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_198_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08031_ _03577_ _03668_ _03579_ _03669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xinput40 la_data_in[4] net40 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_159_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_200_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_174_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_196_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_190_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_171_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09982_ soc.ram_encoder_0.input_buffer\[7\] _04847_ _04248_ _04872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_88_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08933_ _04187_ _00638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_83_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_170_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_85_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_233_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08864_ _04150_ _00606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_229_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_218_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07815_ soc.spi_video_ram_1.write_fifo.fifo_mem\[9\]\[23\] _03460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_111_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3708 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08795_ _04113_ _00574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3719 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_211_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07746_ _02602_ _03390_ _03391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_26_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_225_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_203_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07677_ soc.spi_video_ram_1.write_fifo.fifo_mem\[7\]\[14\] _03323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_26_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_246_1469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_241_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_198_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09416_ _02542_ _04467_ _04471_ _04472_ _00837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_73_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06628_ _02361_ _00160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_90_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_213_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_224_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_209_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09347_ _04424_ _00815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_197_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06559_ _02321_ _00131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_240_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09278_ _03364_ _04375_ _04387_ _00783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_139_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08229_ soc.ram_encoder_0.request_address\[8\] _02505_ _03793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_193_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11240_ _00306_ clknet_leaf_38_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[10\]\[11\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_106_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11171_ _00237_ clknet_leaf_134_wb_clk_i soc.spi_video_ram_1.output_buffer\[19\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_6301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10122_ _04952_ _04967_ _01047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_122_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_231_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_5633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10053_ _04912_ _01034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_103_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4910 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_23_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4921 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_252_wb_clk_i clknet_5_7_0_wb_clk_i clknet_leaf_252_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_4932 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4943 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_1509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5699 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4954 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4965 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4976 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4987 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_217_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4998 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_99_1391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10955_ _00021_ clknet_leaf_255_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[18\]\[9\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_44_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_204_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_186_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_182_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10886_ _05430_ _05431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_147_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_31_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_164_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_73_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_197_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_157_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_200_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_223_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_185_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_157_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11507_ _00573_ clknet_leaf_211_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[23\]\[1\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_32_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_201_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11438_ _00504_ clknet_leaf_72_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[30\]\[19\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_208_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_197_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11369_ _00435_ clknet_leaf_175_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[28\]\[8\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_140_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_10_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_05930_ _01717_ _01823_ _01824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_152_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_230_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05861_ _01563_ soc.cpu.AReg.data\[10\] _01718_ soc.ram_data_out\[10\] _01759_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_26_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_27_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07600_ _03054_ _03246_ _03247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08580_ _02169_ soc.spi_video_ram_1.write_fifo.fifo_mem\[2\]\[24\] _03966_ _03993_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_05792_ _01662_ _01691_ _01693_ _01694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_35_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_207_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07531_ _02919_ _03178_ _03179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_78_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_208_1718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_223_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_228_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07462_ _03054_ _03109_ _03110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_62_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09201_ _01459_ _04346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_06413_ _02230_ _00076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_245_1480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_179_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07393_ soc.spi_video_ram_1.write_fifo.fifo_mem\[14\]\[11\] soc.spi_video_ram_1.write_fifo.fifo_mem\[15\]\[11\]
+ _02613_ _03042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xclkbuf_leaf_56_wb_clk_i clknet_5_13_0_wb_clk_i clknet_leaf_56_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_241_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09132_ _04294_ _04298_ _04299_ _00725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_06344_ _02134_ soc.spi_video_ram_1.write_fifo.fifo_mem\[17\]\[7\] _02182_ _02190_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_104_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09063_ _04261_ _00694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_120_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06275_ soc.spi_video_ram_1.fifo_in_data\[12\] _02145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_175_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08014_ _02685_ _03652_ _02720_ _03653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_50_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_239_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09965_ _04859_ _04848_ _04860_ _00998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_44_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_170_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08916_ soc.spi_video_ram_1.write_fifo.fifo_mem\[22\]\[0\] _02310_ _04178_ _04179_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_103_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09896_ _03765_ _04615_ _04737_ _04808_ _04809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XTAP_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_245_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08847_ _04140_ _00599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_246_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08778_ soc.spi_video_ram_1.write_fifo.fifo_mem\[24\]\[25\] _04069_ _04075_ _04103_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_72_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2804 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2815 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2826 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2837 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07729_ _02655_ _03361_ _03374_ _03375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_2848 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2859 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_3_3_0_wb_clk_i clknet_2_1_0_wb_clk_i clknet_3_3_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_129_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_207_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10740_ soc.spi_video_ram_1.write_fifo.fifo_mem\[31\]\[7\] soc.spi_video_ram_1.fifo_in_data\[7\]
+ _05344_ _05352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_246_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_240_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10671_ _02225_ soc.spi_video_ram_1.write_fifo.fifo_mem\[29\]\[4\] _05310_ _05315_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_129_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12341_ _01369_ clknet_leaf_53_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[8\]\[20\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_139_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_216_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_138_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_1316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12272_ _01300_ clknet_leaf_231_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[31\]\[25\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11223_ _00289_ clknet_leaf_87_wb_clk_i soc.video_generator_1.h_count\[4\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_107_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_194_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6120 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11154_ _00220_ clknet_leaf_165_wb_clk_i soc.ram_encoder_0.output_bits_left\[2\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_218_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6131 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_136_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_6142 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6153 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10105_ soc.ram_data_out\[5\] _04927_ _04954_ _04955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_6164 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_114_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_6175 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11085_ _00151_ clknet_leaf_285_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[13\]\[23\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_95_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_23_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6186 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_49_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_231_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10036_ soc.ram_encoder_0.request_address\[4\] soc.ram_encoder_0.address\[4\] _04900_
+ _04904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_5474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4740 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_49_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4751 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_236_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4762 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4773 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4784 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_149_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4795 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11987_ _01046_ clknet_leaf_158_wb_clk_i soc.ram_data_out\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_1_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_205_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_229_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10938_ soc.spi_video_ram_1.write_fifo.fifo_mem\[8\]\[25\] _04069_ _05430_ _05458_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_56_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_232_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_143_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10869_ _01736_ _05221_ _05412_ _05421_ _01341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_182_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_191_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_185_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06060_ _01946_ _01952_ _01953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_126_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_67_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_154_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_236_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_158_1282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09750_ _04704_ _00939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06962_ _02054_ _02057_ _02623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_234_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_246_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05913_ _01618_ soc.cpu.AReg.data\[13\] _01718_ soc.ram_data_out\[13\] _01808_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_08701_ soc.spi_video_ram_1.write_fifo.fifo_mem\[15\]\[20\] _02343_ _04043_ _04060_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_09681_ _04426_ soc.cpu.PC.REG.data\[6\] _04617_ _04654_ _04655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_171_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_239_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06893_ _02555_ _02558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_228_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08632_ _02159_ soc.spi_video_ram_1.write_fifo.fifo_mem\[30\]\[19\] _04011_ _04021_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_05844_ _01705_ _01742_ _01743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_27_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08563_ _03984_ _00471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_70_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05775_ _01672_ _01676_ _01678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_70_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07514_ _02575_ soc.spi_video_ram_1.write_fifo.fifo_mem\[28\]\[26\] _03161_ _02927_
+ _03162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_74_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08494_ _02145_ soc.spi_video_ram_1.write_fifo.fifo_mem\[28\]\[12\] _03945_ _03948_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_63_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_222_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_1286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07445_ soc.spi_video_ram_1.write_fifo.fifo_mem\[24\]\[27\] soc.spi_video_ram_1.write_fifo.fifo_mem\[25\]\[27\]
+ soc.spi_video_ram_1.write_fifo.fifo_mem\[26\]\[27\] soc.spi_video_ram_1.write_fifo.fifo_mem\[27\]\[27\]
+ _02688_ _02827_ _03094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_168_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_221_1726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07376_ _02922_ soc.spi_video_ram_1.write_fifo.fifo_mem\[17\]\[11\] _03024_ _03025_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_210_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09115_ _02272_ soc.spi_video_ram_1.write_fifo.fifo_mem\[20\]\[27\] _04258_ _04288_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_148_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06327_ _02117_ _02179_ _02180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_191_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09046_ _04247_ _04249_ _00689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06258_ _02133_ _00018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_198_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_150_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06189_ _01542_ _02071_ _02073_ _02075_ _02076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_8_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_132_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_219_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_1279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09948_ _04847_ _04849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_4003 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4014 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_4025 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4036 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09879_ soc.cpu.instruction\[14\] _04741_ _04795_ _04796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_57_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4047 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_3302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_189_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4058 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_218_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4069 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11910_ _00969_ clknet_leaf_128_wb_clk_i soc.cpu.ALU.no vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11841_ _00900_ clknet_leaf_170_wb_clk_i soc.rom_encoder_0.request_data_out\[2\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_73_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1900 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1911 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1922 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_242_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_183_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1933 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11772_ _00833_ clknet_leaf_81_wb_clk_i soc.spi_video_ram_1.read_value\[2\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_57_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1944 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_214_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1955 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1966 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10723_ _05342_ _01274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_53_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1977 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_241_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_198_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1988 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1999 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10654_ _05305_ _01242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_16_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_224_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10585_ net14 _05266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_103_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_202_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12324_ _01352_ clknet_leaf_137_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[8\]\[3\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_177_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_1_wb_clk_i clknet_5_0_0_wb_clk_i clknet_leaf_1_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_177_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12255_ _01283_ clknet_leaf_179_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[31\]\[8\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_126_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_177_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11206_ _00272_ clknet_leaf_26_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[11\]\[16\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12186_ _01214_ net87 soc.gpio_i_stored\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_123_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11137_ _00203_ clknet_leaf_22_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[14\]\[17\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_190_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_235_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_5260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11068_ _00134_ clknet_leaf_208_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[13\]\[6\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_5271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10019_ soc.ram_encoder_0.request_data_out\[12\] soc.ram_encoder_0.data_out\[12\]
+ _04889_ _04895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_49_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_237_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_110_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3880 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_1412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3891 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05560_ soc.spi_video_ram_1.buffer_index\[1\] _01469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_233_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_204_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05491_ soc.spi_video_ram_1.write_fifo.read_pointer\[0\] _01405_ _01406_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_127_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_242_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07230_ _02734_ _02882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_20_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_220_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_165_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_146_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07161_ _02643_ _02815_ _02816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_30_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06112_ soc.video_generator_1.h_count\[2\] _01902_ _02005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_07092_ soc.spi_video_ram_1.write_fifo.fifo_mem\[8\]\[3\] soc.spi_video_ram_1.write_fifo.fifo_mem\[9\]\[3\]
+ soc.spi_video_ram_1.write_fifo.fifo_mem\[10\]\[3\] soc.spi_video_ram_1.write_fifo.fifo_mem\[11\]\[3\]
+ _02713_ _02714_ _02749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_246_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06043_ _01928_ _01929_ _01935_ _01936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_132_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09802_ _02459_ _04731_ _04733_ _04734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_134_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07994_ _03627_ _03629_ _03631_ _03633_ _02568_ _03634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_68_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09733_ _04677_ _04693_ _04694_ _01381_ _00932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_06945_ _01391_ _02606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_60_1747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_214_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_83_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09664_ _04642_ soc.rom_encoder_0.request_address\[1\] _04632_ _04643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06876_ _02544_ _00225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_227_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05827_ _01711_ _01726_ _01727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_08615_ _04012_ _00495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_83_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09595_ soc.rom_encoder_0.input_buffer\[6\] _04598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_167_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_71_wb_clk_i clknet_5_9_0_wb_clk_i clknet_leaf_71_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_224_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_208_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05758_ _01635_ _01647_ _01649_ _01662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_39_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08546_ _03975_ _00463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_211_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_223_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08477_ _02128_ soc.spi_video_ram_1.write_fifo.fifo_mem\[28\]\[4\] _03934_ _03939_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_05689_ _01558_ soc.cpu.ALU.x\[1\] _01596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_51_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07428_ _02597_ soc.spi_video_ram_1.write_fifo.fifo_mem\[6\]\[27\] _02690_ _03077_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_17_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_196_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_109_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_149_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07359_ _03005_ _03006_ _03008_ _02908_ _02581_ _03009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_137_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_137_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xcaravel_hack_soc_104 io_oeb[21] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xcaravel_hack_soc_115 io_out[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_10370_ _05126_ _01137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_100_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xcaravel_hack_soc_126 irq[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xcaravel_hack_soc_137 la_data_out[9] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xcaravel_hack_soc_148 la_data_out[20] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xcaravel_hack_soc_159 la_data_out[32] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_09029_ _03338_ _04224_ _04238_ _00683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_3_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_151_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_1731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12040_ _01099_ clknet_leaf_274_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[5\]\[28\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_156_1753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_5_24_0_wb_clk_i clknet_4_12_0_wb_clk_i clknet_5_24_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_46_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_191_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_232_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_1_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_150_1352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3110 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_219_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3121 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3132 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_185_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3143 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_233_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3154 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_34_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3165 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3176 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3187 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11824_ _00883_ clknet_leaf_96_wb_clk_i soc.rom_encoder_0.input_bits_left\[3\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1730 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_215_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1752 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1763 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11755_ _00816_ clknet_leaf_279_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[4\]\[28\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1785 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1796 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_202_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10706_ _02258_ soc.spi_video_ram_1.write_fifo.fifo_mem\[29\]\[20\] _05321_ _05334_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_187_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11686_ _00747_ clknet_leaf_142_wb_clk_i soc.spi_video_ram_1.fifo_in_data\[4\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10637_ soc.spi_video_ram_1.write_fifo.fifo_mem\[19\]\[17\] soc.spi_video_ram_1.fifo_in_address\[1\]
+ _05289_ _05297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_70_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10568_ _05173_ _05254_ _05255_ _01206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_220_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12307_ _01335_ clknet_leaf_144_wb_clk_i soc.ram_encoder_0.data_out\[2\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_143_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_196_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10499_ soc.cpu.PC.REG.data\[13\] _05212_ _05213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_83_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_216_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_155_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12238_ _01266_ clknet_leaf_49_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[29\]\[20\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_130_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12169_ _01197_ clknet_leaf_154_wb_clk_i soc.ram_encoder_0.address\[14\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_25_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_211_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput5 io_in[16] net5 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyd_1
X_06730_ soc.spi_video_ram_1.write_fifo.fifo_mem\[14\]\[17\] _02337_ _02412_ _02421_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_211_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5090 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_209_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_188_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_06661_ _02378_ _00176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_227_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08400_ soc.spi_video_ram_1.write_fifo.fifo_mem\[26\]\[28\] _02353_ _03865_ _03896_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_05612_ _01516_ _01517_ _01519_ _01520_ _01521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_206_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_149_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09380_ soc.spi_video_ram_1.state_sram_clk_counter\[7\] _04445_ _04447_ _00825_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_209_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06592_ soc.spi_video_ram_1.write_fifo.fifo_mem\[13\]\[18\] _02339_ _02328_ _02340_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_178_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_196_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08331_ _03858_ _00365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05543_ soc.ram_encoder_0.initialized soc.rom_encoder_0.initialized soc.spi_video_ram_1.initialized
+ _01453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_33_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_205_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08262_ _03815_ _03818_ _03819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_60_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05474_ _01388_ _01389_ _01390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_127_1387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_221_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_178_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07213_ soc.spi_video_ram_1.write_fifo.fifo_mem\[0\]\[8\] soc.spi_video_ram_1.write_fifo.fifo_mem\[1\]\[8\]
+ soc.spi_video_ram_1.write_fifo.fifo_mem\[2\]\[8\] soc.spi_video_ram_1.write_fifo.fifo_mem\[3\]\[8\]
+ _02591_ _02593_ _02865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_192_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08193_ _03762_ _00323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_119_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_146_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07144_ _02793_ _02795_ _02797_ _02799_ _02568_ _02800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_118_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07075_ _02674_ _00830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_161_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06026_ _01876_ _01917_ _01919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_161_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_236_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_5_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07977_ soc.spi_video_ram_1.write_fifo.fifo_mem\[8\]\[18\] soc.spi_video_ram_1.write_fifo.fifo_mem\[9\]\[18\]
+ soc.spi_video_ram_1.write_fifo.fifo_mem\[10\]\[18\] soc.spi_video_ram_1.write_fifo.fifo_mem\[11\]\[18\]
+ _02701_ _02737_ _03617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_102_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09716_ _04679_ _04680_ _03778_ soc.ram_encoder_0.output_buffer\[16\] _04681_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_5_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06928_ _02588_ _02589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_99_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_215_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09647_ _04617_ _04632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_16_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06859_ _01822_ _01825_ _02529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_28_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_231_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09578_ net5 _04586_ _04553_ _04587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_145_1410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_227_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08529_ _03965_ _03966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_169_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_277_wb_clk_i clknet_5_4_0_wb_clk_i clknet_leaf_277_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_11540_ _00606_ clknet_leaf_179_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[25\]\[5\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_204_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11471_ _00537_ clknet_leaf_284_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[15\]\[23\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_51_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10422_ _02272_ soc.spi_video_ram_1.write_fifo.fifo_mem\[6\]\[27\] _05123_ _05153_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_104_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_193_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_87_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10353_ _01767_ _05104_ _05116_ _01130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_109_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10284_ soc.rom_loader.current_address\[1\] _05069_ _05070_ _05073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_2_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_1403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12023_ _01082_ clknet_leaf_38_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[5\]\[11\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_105_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_215_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_78_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_185_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_234_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_221_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_178_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11807_ _00867_ clknet_leaf_288_wb_clk_i soc.spi_video_ram_1.fifo_in_address\[10\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_128_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_1505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11738_ _00799_ clknet_leaf_39_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[4\]\[11\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_203_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_187_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11669_ _00730_ clknet_leaf_64_wb_clk_i soc.spi_video_ram_1.state_counter\[8\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_70_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_190_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_190_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_183_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_115_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_44_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_233_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07900_ _03047_ soc.spi_video_ram_1.write_fifo.fifo_mem\[14\]\[21\] _03542_ _02652_
+ _03543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_9_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08880_ soc.spi_video_ram_1.write_fifo.fifo_mem\[25\]\[13\] _04050_ _04155_ _04159_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_44_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07831_ soc.spi_video_ram_1.output_buffer\[8\] _02882_ _03473_ _03475_ _03476_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_99_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_244_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07762_ _02952_ _03403_ _03406_ _03407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_238_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09501_ _04535_ _00859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06713_ soc.spi_video_ram_1.fifo_in_data\[10\] _02411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_07693_ _02612_ _03338_ _03339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_77_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_168_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_213_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09432_ soc.rom_encoder_0.request_address\[10\] _02520_ _04460_ soc.rom_encoder_0.output_buffer\[7\]
+ _04484_ _04485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_06644_ _02143_ soc.spi_video_ram_1.write_fifo.fifo_mem\[12\]\[11\] _02368_ _02370_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_92_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_80_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_197_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_146_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_06575_ soc.spi_video_ram_1.write_fifo.fifo_mem\[13\]\[11\] _02240_ _02328_ _02330_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_09363_ _04435_ _04436_ _00819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_181_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_33_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08314_ _02155_ soc.spi_video_ram_1.write_fifo.fifo_mem\[1\]\[17\] _03842_ _03850_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_05526_ _01437_ _01424_ _01438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_244_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_162_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09294_ _04397_ _00789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_123_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_205_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_10 net76 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08245_ soc.ram_encoder_0.request_address\[12\] _02505_ _03805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_193_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_197_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08176_ _02161_ soc.spi_video_ram_1.write_fifo.fifo_mem\[10\]\[20\] _03731_ _03754_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_105_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_238_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_179_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07127_ _02573_ _02783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
X_07058_ _02712_ _02717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XTAP_6505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06009_ soc.display_clks_before_active\[0\] _01842_ _01902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_121_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_6538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5804 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5815 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_47_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5826 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_212_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5837 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5848 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5859 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_134_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_228_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_186_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10971_ _00037_ clknet_leaf_234_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[18\]\[25\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_95_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_216_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_203_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_223_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11523_ _00589_ clknet_leaf_29_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[23\]\[17\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_183_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_172_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11454_ _00520_ clknet_leaf_202_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[15\]\[6\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_125_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10405_ _05144_ _01154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_11385_ _00451_ clknet_leaf_300_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[28\]\[24\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_152_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_125_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10336_ _01632_ _05103_ _05107_ _01122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_112_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10267_ _02274_ soc.spi_video_ram_1.write_fifo.fifo_mem\[5\]\[28\] _05041_ _05062_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_79_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_238_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_12006_ _01065_ clknet_leaf_113_wb_clk_i soc.hack_clock_0.counter\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_152_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_61_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10198_ soc.hack_clock_0.counter\[4\] _05022_ _05024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_234_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_43_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_226_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_228_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xclkbuf_leaf_199_wb_clk_i clknet_5_18_0_wb_clk_i clknet_leaf_199_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_98_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_179_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xclkbuf_leaf_128_wb_clk_i clknet_5_13_0_wb_clk_i clknet_leaf_128_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_2080 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2091 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_163_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06360_ _02198_ _00055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_188_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06291_ _02155_ soc.spi_video_ram_1.write_fifo.fifo_mem\[18\]\[17\] _02141_ _02156_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_50_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08030_ soc.spi_video_ram_1.write_fifo.fifo_mem\[28\]\[16\] soc.spi_video_ram_1.write_fifo.fifo_mem\[29\]\[16\]
+ soc.spi_video_ram_1.write_fifo.fifo_mem\[30\]\[16\] soc.spi_video_ram_1.write_fifo.fifo_mem\[31\]\[16\]
+ _02726_ _03041_ _03668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
Xinput30 la_data_in[20] net30 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput41 la_data_in[5] net41 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_239_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_4_5_0_wb_clk_i clknet_3_2_0_wb_clk_i clknet_4_5_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_85_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_192_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09981_ soc.ram_encoder_0.input_buffer\[11\] _04871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_171_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_100_1390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08932_ soc.spi_video_ram_1.write_fifo.fifo_mem\[22\]\[8\] _02407_ _04178_ _04187_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_112_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_213_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08863_ soc.spi_video_ram_1.write_fifo.fifo_mem\[25\]\[5\] _02401_ _04144_ _04150_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_135_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07814_ _02704_ soc.spi_video_ram_1.write_fifo.fifo_mem\[11\]\[23\] _02593_ _03459_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_111_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3709 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08794_ _02124_ soc.spi_video_ram_1.write_fifo.fifo_mem\[23\]\[2\] _04110_ _04113_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_245_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07745_ _03385_ _03386_ _03389_ _02952_ _03390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_84_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_168_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07676_ _02574_ soc.spi_video_ram_1.write_fifo.fifo_mem\[4\]\[14\] _03321_ _02740_
+ _03322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_38_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_240_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09415_ soc.rom_encoder_0.output_buffer\[7\] _02541_ _04472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_53_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06627_ _02126_ soc.spi_video_ram_1.write_fifo.fifo_mem\[12\]\[3\] _02357_ _02361_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_09346_ _02272_ soc.spi_video_ram_1.write_fifo.fifo_mem\[4\]\[27\] _04394_ _04424_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06558_ soc.spi_video_ram_1.write_fifo.fifo_mem\[13\]\[3\] _02223_ _02317_ _02321_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_224_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05509_ soc.spi_video_ram_1.state_sram_clk_counter\[3\] soc.spi_video_ram_1.state_sram_clk_counter\[2\]
+ _01388_ _01416_ _01424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_225_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09277_ _04067_ _04360_ _04387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06489_ _02124_ soc.spi_video_ram_1.write_fifo.fifo_mem\[0\]\[2\] _02279_ _02282_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_166_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08228_ _02556_ _03791_ _03792_ _00328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_154_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_140_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08159_ _03745_ _00306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_101_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_162_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_218_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_162_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11170_ _00236_ clknet_leaf_136_wb_clk_i soc.spi_video_ram_1.output_buffer\[20\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_161_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_175_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10121_ soc.ram_data_out\[9\] _04927_ _04966_ _04967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_6324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_216_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_231_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_5601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10052_ soc.ram_encoder_0.request_address\[12\] soc.ram_encoder_0.address\[12\] _04879_
+ _04912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4900 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_130_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_196_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_88_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_236_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4911 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4922 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_130_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4933 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_180_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_208_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4944 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4955 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4966 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_169_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_235_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4977 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_169_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4988 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4999 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_17_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_292_wb_clk_i clknet_5_5_0_wb_clk_i clknet_leaf_292_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_91_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_232_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_229_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10954_ _00020_ clknet_leaf_219_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[18\]\[8\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_56_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_221_wb_clk_i clknet_5_23_0_wb_clk_i clknet_leaf_221_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_95_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10885_ _05429_ _05430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_108_1319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_231_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_106_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_106_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_185_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11506_ _00572_ clknet_5_22_0_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[23\]\[0\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_240_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11437_ _00503_ clknet_leaf_73_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[30\]\[18\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_153_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_193_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11368_ _00434_ clknet_leaf_186_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[28\]\[7\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_153_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10319_ _05070_ _05095_ _05096_ _01115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_154_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11299_ _00365_ clknet_leaf_229_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[1\]\[25\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_112_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_239_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_224_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_152_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05860_ _01557_ _01757_ _01758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_227_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_309_wb_clk_i clknet_5_1_0_wb_clk_i clknet_leaf_309_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_94_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05791_ _01677_ _01692_ _01693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_47_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07530_ soc.spi_video_ram_1.write_fifo.fifo_mem\[5\]\[26\] _03178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_19_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_78_1476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_222_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07461_ soc.spi_video_ram_1.write_fifo.fifo_mem\[23\]\[12\] _03109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_35_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_17_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06412_ soc.spi_video_ram_1.write_fifo.fifo_mem\[16\]\[6\] _02229_ _02217_ _02230_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_91_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09200_ _00011_ _01666_ _04345_ _00747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_210_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07392_ _02958_ _03041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_72_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_206_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06343_ _02189_ _00047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09131_ soc.spi_video_ram_1.state_counter\[3\] _04296_ _04299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_33_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_31_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_191_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_147_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09062_ _02219_ soc.spi_video_ram_1.write_fifo.fifo_mem\[20\]\[1\] _04259_ _04261_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_198_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06274_ _02144_ _00023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xclkbuf_leaf_96_wb_clk_i clknet_5_11_0_wb_clk_i clknet_leaf_96_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_50_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_200_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08013_ soc.spi_video_ram_1.write_fifo.fifo_mem\[20\]\[17\] soc.spi_video_ram_1.write_fifo.fifo_mem\[21\]\[17\]
+ soc.spi_video_ram_1.write_fifo.fifo_mem\[22\]\[17\] soc.spi_video_ram_1.write_fifo.fifo_mem\[23\]\[17\]
+ _02717_ _02682_ _03652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_85_1414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_25_wb_clk_i clknet_5_8_0_wb_clk_i clknet_leaf_25_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_190_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_235_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09964_ soc.ram_encoder_0.input_buffer\[1\] _04849_ _04248_ _04860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_104_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_217_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08915_ _04177_ _04178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_09895_ _02437_ _04807_ _04808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_218_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08846_ _02175_ soc.spi_video_ram_1.write_fifo.fifo_mem\[23\]\[27\] _04109_ _04140_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_246_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_217_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08777_ _04102_ _00567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2805 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_175_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05989_ _01853_ soc.video_generator_1.v_count\[0\] _01850_ soc.boot_loading_offset\[0\]
+ _01882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_26_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2816 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2827 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_214_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07728_ _02585_ _03367_ _03373_ _03374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_2838 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2849 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_241_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_198_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_183_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07659_ _03288_ _03295_ _03304_ _03305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_213_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_246_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_224_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10670_ _05314_ _01249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_16_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_55_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_70_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09329_ _04415_ _00806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_70_1749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_194_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12340_ _01368_ clknet_leaf_31_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[8\]\[19\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_193_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12271_ _01299_ clknet_leaf_299_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[31\]\[24\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_5_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_209_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_182_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11222_ _00288_ clknet_leaf_87_wb_clk_i soc.video_generator_1.h_count\[3\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_120_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_190_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6110 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11153_ _00219_ clknet_leaf_166_wb_clk_i soc.ram_encoder_0.output_bits_left\[3\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_122_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6121 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6132 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6143 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10104_ _04851_ _04947_ _04948_ _04953_ _04954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_6154 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11084_ _00150_ clknet_leaf_267_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[13\]\[22\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_6165 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_6176 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_88_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6187 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_49_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_237_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10035_ _04903_ _01025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_5464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4730 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_209_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4741 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4752 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_4763 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4774 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4785 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4796 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11986_ _01045_ clknet_leaf_144_wb_clk_i soc.ram_data_out\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_204_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_182_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10937_ _05457_ _01373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_95_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_189_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10868_ soc.ram_encoder_0.data_out\[8\] _05421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_158_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_160_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_223_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10799_ _02227_ soc.spi_video_ram_1.write_fifo.fifo_mem\[7\]\[5\] _05378_ _05384_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_34_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_184_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_199_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_158_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_185_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_201_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_172_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_214_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06961_ _02606_ _02621_ _02622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_79_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_230_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08700_ _04059_ _00533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05912_ _01702_ _01806_ _01807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_45_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09680_ _04639_ soc.rom_loader.current_address\[6\] _04654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_06892_ soc.ram_encoder_0.request_address\[3\] _02506_ _02557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_67_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_143_wb_clk_i clknet_5_24_0_wb_clk_i clknet_leaf_143_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_82_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08631_ _04020_ _00503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05843_ _01717_ _01741_ _01742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_95_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08562_ _02151_ soc.spi_video_ram_1.write_fifo.fifo_mem\[2\]\[15\] _03978_ _03984_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_05774_ _01672_ _01676_ _01677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_223_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07513_ _02903_ _03160_ _03161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_93_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_50_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08493_ _03947_ _00438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_62_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07444_ _02719_ _03087_ _03092_ _03093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_149_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_211_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_241_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07375_ _02741_ _03024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_176_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09114_ _04287_ _00719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_13_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06326_ soc.spi_video_ram_1.write_fifo.write_pointer\[1\] _01444_ _02179_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_149_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_175_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06257_ _02132_ soc.spi_video_ram_1.write_fifo.fifo_mem\[18\]\[6\] _02120_ _02133_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_09045_ soc.spi_video_ram_1.write_fifo.read_pointer\[1\] _04246_ _04248_ _04249_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_191_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_209_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_191_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_239_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06188_ _01519_ _01543_ _01545_ _01523_ _02074_ _02075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
Xclkbuf_5_14_0_wb_clk_i clknet_4_7_0_wb_clk_i clknet_5_14_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_89_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09947_ _04847_ _04848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_8_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_63_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4004 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_219_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4015 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09878_ _04607_ _04743_ _04739_ _04794_ _04795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_4026 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4037 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_213_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4048 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4059 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08829_ _04131_ _00590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11840_ _00899_ clknet_5_11_0_wb_clk_i soc.rom_encoder_0.request_data_out\[1\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1901 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1923 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_199_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11771_ _00832_ clknet_leaf_82_wb_clk_i soc.spi_video_ram_1.read_value\[1\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1934 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1945 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1956 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10722_ _02274_ soc.spi_video_ram_1.write_fifo.fifo_mem\[29\]\[28\] _05321_ _05342_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_1967 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1978 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1989 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_201_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10653_ soc.spi_video_ram_1.write_fifo.fifo_mem\[19\]\[25\] _04069_ _05277_ _05305_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_16_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_220_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10584_ _01652_ _05261_ _05265_ _01212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_16_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_177_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12323_ _01351_ clknet_leaf_137_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[8\]\[2\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_182_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_107_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12254_ _01282_ clknet_leaf_193_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[31\]\[7\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_194_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11205_ _00271_ clknet_leaf_8_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[11\]\[15\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12185_ _01213_ net86 soc.gpio_i_stored\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_69_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_218_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_1478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_150_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11136_ _00202_ clknet_leaf_20_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[14\]\[16\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_96_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_231_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_133_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11067_ _00133_ clknet_leaf_219_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[13\]\[5\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_5261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_7_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_49_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10018_ _04894_ _01017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_77_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_236_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_110_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3870 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3881 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_205_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3892 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11969_ _01028_ clknet_leaf_183_wb_clk_i soc.ram_encoder_0.request_address\[6\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_229_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_244_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_232_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_166_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05490_ soc.spi_video_ram_1.write_fifo.write_pointer\[0\] _01405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_53_1722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07160_ soc.spi_video_ram_1.write_fifo.fifo_mem\[16\]\[5\] soc.spi_video_ram_1.write_fifo.fifo_mem\[17\]\[5\]
+ soc.spi_video_ram_1.write_fifo.fifo_mem\[18\]\[5\] soc.spi_video_ram_1.write_fifo.fifo_mem\[19\]\[5\]
+ _02645_ _02647_ _02815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_185_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_160_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_121_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06111_ _01924_ _01984_ _02004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_9_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07091_ _02736_ _02738_ _02747_ _02720_ _02748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_121_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_246_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06042_ soc.boot_loading_offset\[4\] _01934_ _01935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_236_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09801_ _02459_ _04732_ _04733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_119_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07993_ _02685_ _03632_ _03579_ _03633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_140_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09732_ net61 _04677_ _04694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_171_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06944_ _02568_ _02604_ _02605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_67_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_228_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09663_ soc.cpu.PC.REG.data\[1\] soc.rom_loader.current_address\[1\] _04639_ _04642_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06875_ soc.rom_encoder_0.output_buffer\[4\] _02542_ _02543_ soc.rom_encoder_0.request_address\[3\]
+ _02544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_54_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08614_ _02140_ soc.spi_video_ram_1.write_fifo.fifo_mem\[30\]\[10\] _04011_ _04012_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_05826_ _01696_ _01710_ _01726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09594_ _04596_ _04585_ _04597_ _00890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_70_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08545_ _02134_ soc.spi_video_ram_1.write_fifo.fifo_mem\[2\]\[7\] _03967_ _03975_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_05757_ _01656_ _01660_ _01661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_184_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08476_ _03938_ _00430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_126_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05688_ _01594_ _01595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_208_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07427_ _02941_ soc.spi_video_ram_1.write_fifo.fifo_mem\[7\]\[27\] _03076_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_7_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_40_wb_clk_i clknet_5_3_0_wb_clk_i clknet_leaf_40_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_104_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_210_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_164_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07358_ _02695_ soc.spi_video_ram_1.write_fifo.fifo_mem\[28\]\[28\] _03007_ _03008_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_221_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xcaravel_hack_soc_105 io_oeb[27] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_06309_ _02167_ soc.spi_video_ram_1.write_fifo.fifo_mem\[18\]\[23\] _02119_ _02168_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xcaravel_hack_soc_116 io_out[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_152_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xcaravel_hack_soc_127 irq[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_07289_ _02696_ soc.spi_video_ram_1.write_fifo.fifo_mem\[7\]\[10\] _02939_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_136_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xcaravel_hack_soc_138 la_data_out[10] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_09028_ _04067_ _04225_ _04238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xcaravel_hack_soc_149 la_data_out[21] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_163_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_137_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_219_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_172_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_172_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3100 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_218_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3111 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3122 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3133 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_111_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3144 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_3155 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_234_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3166 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3177 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11823_ _00882_ clknet_leaf_96_wb_clk_i soc.rom_encoder_0.input_bits_left\[2\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1720 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_57_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_233_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_183_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1731 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_214_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_26_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1742 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_183_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1753 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1764 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11754_ _00815_ clknet_5_6_0_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[4\]\[27\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_226_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1775 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_230_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_198_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1786 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1797 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10705_ _05333_ _01265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_109_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11685_ _00746_ clknet_leaf_132_wb_clk_i soc.spi_video_ram_1.fifo_in_data\[3\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_224_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_186_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10636_ _05296_ _01233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_167_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_161_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10567_ net19 _05255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_6_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_155_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12306_ _01334_ clknet_leaf_144_wb_clk_i soc.ram_encoder_0.data_out\[1\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_115_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10498_ soc.cpu.PC.REG.data\[11\] soc.cpu.PC.REG.data\[12\] _05206_ _05212_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_12237_ _01265_ clknet_leaf_71_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[29\]\[19\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_237_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_1245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12168_ _01196_ clknet_leaf_152_wb_clk_i soc.ram_encoder_0.address\[13\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_151_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_190_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11119_ _00185_ clknet_leaf_281_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[12\]\[28\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_46_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12099_ _01127_ net86 soc.cpu.ALU.x\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_232_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput6 io_in[17] net6 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XTAP_5080 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_110_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_237_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5091 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06660_ _02159_ soc.spi_video_ram_1.write_fifo.fifo_mem\[12\]\[19\] _02368_ _02378_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_4390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_52_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05611_ soc.spi_video_ram_1.output_buffer\[10\] soc.spi_video_ram_1.output_buffer\[11\]
+ _01468_ _01520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06591_ soc.spi_video_ram_1.fifo_in_address\[2\] _02339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_51_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_233_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08330_ _02171_ soc.spi_video_ram_1.write_fifo.fifo_mem\[1\]\[25\] _03830_ _03858_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_05542_ soc.rom_encoder_0.write_enable net18 net13 net37 _01452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or4_2
XFILLER_178_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_166_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_209_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08261_ _03816_ _02510_ _03788_ soc.ram_encoder_0.request_data_out\[8\] _03817_ _03818_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_05473_ soc.spi_video_ram_1.state_sram_clk_counter\[3\] soc.spi_video_ram_1.state_sram_clk_counter\[2\]
+ _01389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_220_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07212_ _02571_ _02863_ _02586_ _02864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_14_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08192_ _02177_ soc.spi_video_ram_1.write_fifo.fifo_mem\[10\]\[28\] _03731_ _03762_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_9_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07143_ _02768_ _02798_ _02799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_101_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07074_ _02677_ _02606_ _02711_ _02732_ _02733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_145_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06025_ _01876_ _01917_ _01918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_86_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_43_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07976_ _01539_ _02882_ _03596_ _03616_ _00252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_45_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_214_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09715_ _02482_ _02499_ _04680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_142_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06927_ _02581_ _02588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_19_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09646_ _04631_ _00908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_216_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06858_ soc.cpu.AReg.data\[15\] _02528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_186_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05809_ _01704_ _01709_ _01710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09577_ _04584_ _04586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06789_ net65 _02453_ _02468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_215_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_145_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08528_ _02114_ _02276_ _03965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_212_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_243_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08459_ soc.spi_video_ram_1.write_fifo.fifo_mem\[27\]\[26\] _03927_ _03898_ _03928_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_184_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_196_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_225_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_211_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11470_ _00536_ clknet_leaf_268_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[15\]\[22\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_184_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_177_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10421_ _05152_ _01162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_109_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_246_wb_clk_i clknet_5_17_0_wb_clk_i clknet_leaf_246_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_100_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10352_ soc.cpu.ALU.x\[10\] _05109_ _05116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_192_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_151_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10283_ _05069_ _05071_ _05072_ _01103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_152_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_65_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12022_ _01081_ clknet_leaf_15_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[5\]\[10\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_133_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_191_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_232_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_219_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xclkbuf_5_7_0_wb_clk_i clknet_4_3_0_wb_clk_i clknet_5_7_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_46_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_185_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_215_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11806_ _00866_ clknet_leaf_288_wb_clk_i soc.spi_video_ram_1.fifo_in_address\[9\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_199_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11737_ _00798_ clknet_leaf_15_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[4\]\[10\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_72_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_202_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_124_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11668_ _00729_ clknet_leaf_66_wb_clk_i soc.spi_video_ram_1.state_counter\[7\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_70_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10619_ _05287_ _01225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_204_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11599_ _00665_ clknet_leaf_248_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[21\]\[6\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_157_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_128_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_183_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_196_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_182_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_124_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_29_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_1556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07830_ _03474_ _02625_ _02882_ _03475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_81_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07761_ _02784_ soc.spi_video_ram_1.write_fifo.fifo_mem\[14\]\[15\] _03405_ _02647_
+ _03406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_37_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09500_ _02254_ soc.cpu.AReg.data\[2\] _04339_ _04535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06712_ _02410_ _00195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07692_ soc.spi_video_ram_1.write_fifo.fifo_mem\[21\]\[24\] _03338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_1601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09431_ soc.rom_encoder_0.request_data_out\[3\] _03767_ _04484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_37_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06643_ _02369_ _00167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_164_1319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09362_ soc.spi_video_ram_1.state_sram_clk_counter\[1\] _04432_ _04433_ _04436_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06574_ _02329_ _00138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_146_1753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08313_ _03849_ _00356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05525_ soc.spi_video_ram_1.current_state\[1\] _01437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_127_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09293_ _02219_ soc.spi_video_ram_1.write_fifo.fifo_mem\[4\]\[1\] _04395_ _04397_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_20_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_11 net83 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_221_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_178_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08244_ _02558_ _03803_ _03804_ _00332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_192_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_222_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08175_ _03753_ _00314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_140_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07126_ soc.spi_video_ram_1.write_fifo.fifo_mem\[8\]\[4\] soc.spi_video_ram_1.write_fifo.fifo_mem\[9\]\[4\]
+ soc.spi_video_ram_1.write_fifo.fifo_mem\[10\]\[4\] soc.spi_video_ram_1.write_fifo.fifo_mem\[11\]\[4\]
+ _02713_ _02714_ _02782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_49_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07057_ _02678_ _02715_ _02716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_6506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06008_ soc.video_generator_1.h_count\[3\] _01842_ _01901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_47_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_5805 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_138_1281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_5816 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5827 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_173_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5838 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_87_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5849 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_29_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07959_ soc.spi_video_ram_1.write_fifo.fifo_mem\[12\]\[19\] soc.spi_video_ram_1.write_fifo.fifo_mem\[13\]\[19\]
+ soc.spi_video_ram_1.write_fifo.fifo_mem\[14\]\[19\] soc.spi_video_ram_1.write_fifo.fifo_mem\[15\]\[19\]
+ _02701_ _02737_ _03600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_46_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10970_ _00036_ clknet_leaf_301_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[18\]\[24\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_21_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_210_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09629_ soc.rom_encoder_0.data_out\[2\] soc.rom_encoder_0.request_data_out\[2\] _04621_
+ _04623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_95_1438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_244_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_239_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_197_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11522_ _00588_ clknet_leaf_29_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[23\]\[16\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_240_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_141_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_201_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11453_ _00519_ clknet_leaf_222_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[15\]\[5\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_201_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10404_ _02254_ soc.spi_video_ram_1.write_fifo.fifo_mem\[6\]\[18\] _05135_ _05144_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_11384_ _00450_ clknet_leaf_290_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[28\]\[23\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_139_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_164_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_217_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10335_ soc.cpu.ALU.x\[2\] _05104_ _05107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_238_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_152_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10266_ _05061_ _01098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_87_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_65_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_12005_ _01064_ clknet_leaf_115_wb_clk_i soc.hack_clock_0.counter\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_120_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10197_ _05017_ _05022_ _05023_ _01067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_121_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_238_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_35_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_234_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_185_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_62_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2070 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2081 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_50_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2092 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_203_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_175_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_226_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_168_wb_clk_i clknet_5_30_0_wb_clk_i clknet_leaf_168_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_06290_ soc.spi_video_ram_1.fifo_in_address\[1\] _02155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_174_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput20 la_data_in[11] net20 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput31 la_data_in[21] net31 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_190_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xinput42 la_data_in[6] net42 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_162_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09980_ _04869_ _04849_ _04870_ _01003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_66_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08931_ _04186_ _00637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_217_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08862_ _04149_ _00605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_69_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07813_ _03047_ soc.spi_video_ram_1.write_fifo.fifo_mem\[10\]\[23\] _03458_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_111_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08793_ _04112_ _00573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_244_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07744_ _02784_ soc.spi_video_ram_1.write_fifo.fifo_mem\[20\]\[15\] _03388_ _03024_
+ _03389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_26_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_77_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_226_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07675_ _02902_ _03320_ _03321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_16_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09414_ _04469_ _04470_ _04471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_52_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06626_ _02360_ _00159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_197_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_201_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09345_ _04423_ _00814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06557_ _02320_ _00130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_244_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_205_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05508_ soc.spi_video_ram_1.state_sram_clk_counter\[6\] soc.spi_video_ram_1.state_sram_clk_counter\[5\]
+ soc.spi_video_ram_1.state_sram_clk_counter\[4\] _01422_ _01423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
X_09276_ _03460_ _04375_ _04386_ _00782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_193_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06488_ _02281_ _00100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_194_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08227_ soc.ram_encoder_0.output_buffer\[8\] _02563_ _03792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_105_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08158_ _02143_ soc.spi_video_ram_1.write_fifo.fifo_mem\[10\]\[11\] _03743_ _03745_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_146_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07109_ _02571_ _02765_ _02586_ _02766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08089_ soc.spi_video_ram_1.write_fifo.fifo_mem\[11\]\[22\] _02262_ _03679_ _03704_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_84_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10120_ _04859_ _04947_ _04948_ _04965_ _04966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_122_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_192_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10051_ _04911_ _01033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_27_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4901 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4912 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4923 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4934 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4945 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4956 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4967 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_4978 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_91_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4989 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10953_ _00019_ clknet_leaf_194_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[18\]\[7\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_189_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_216_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10884_ _02214_ _03729_ _05429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_232_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_223_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_73_1555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_160_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xclkbuf_leaf_261_wb_clk_i clknet_5_7_0_wb_clk_i clknet_leaf_261_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XPHY_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_185_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11505_ _00571_ clknet_leaf_297_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[24\]\[28\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_172_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_32_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11436_ _00502_ clknet_leaf_76_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[30\]\[17\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_171_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11367_ _00433_ clknet_leaf_208_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[28\]\[6\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_67_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10318_ soc.rom_loader.current_address\[12\] _05094_ _05096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_11298_ _00364_ clknet_leaf_296_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[1\]\[24\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_136_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_171_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10249_ _02256_ soc.spi_video_ram_1.write_fifo.fifo_mem\[5\]\[19\] _05041_ _05053_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_26_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_234_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_226_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_239_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_187_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05790_ _01656_ _01660_ _01672_ _01676_ _01692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_94_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_240_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_228_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_169_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_208_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07460_ soc.spi_video_ram_1.write_fifo.fifo_mem\[16\]\[12\] soc.spi_video_ram_1.write_fifo.fifo_mem\[17\]\[12\]
+ soc.spi_video_ram_1.write_fifo.fifo_mem\[18\]\[12\] soc.spi_video_ram_1.write_fifo.fifo_mem\[19\]\[12\]
+ _02903_ _02904_ _03108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_126_1409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06411_ soc.spi_video_ram_1.fifo_in_data\[6\] _02229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_50_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07391_ _02620_ _03032_ _03039_ _03040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_245_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_188_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09130_ soc.spi_video_ram_1.state_counter\[3\] _04296_ _04298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_06342_ _02132_ soc.spi_video_ram_1.write_fifo.fifo_mem\[17\]\[6\] _02182_ _02189_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_202_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09061_ _04260_ _00693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_120_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06273_ _02143_ soc.spi_video_ram_1.write_fifo.fifo_mem\[18\]\[11\] _02141_ _02144_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_191_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08012_ _02678_ _03650_ _03651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_163_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_128_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09963_ soc.ram_encoder_0.input_buffer\[5\] _04859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_103_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xclkbuf_leaf_65_wb_clk_i clknet_5_11_0_wb_clk_i clknet_leaf_65_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_08914_ _04176_ _04177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_213_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09894_ _02433_ _04730_ _02450_ _04807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08845_ _03151_ _04124_ _04139_ _00598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_245_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08776_ soc.spi_video_ram_1.write_fifo.fifo_mem\[24\]\[24\] _04067_ _04075_ _04102_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_3529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05988_ soc.boot_loading_offset\[3\] _01881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_22_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2806 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2817 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07727_ _02900_ _03370_ _03372_ _03373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_2828 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_232_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2839 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_129_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_246_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07658_ _02642_ _03296_ _03303_ _02585_ _03304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_246_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_246_1279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_214_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_186_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06609_ _02349_ _00153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07589_ _02693_ _03232_ _03235_ _02901_ _03236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_139_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09328_ _02254_ soc.spi_video_ram_1.write_fifo.fifo_mem\[4\]\[18\] _04406_ _04415_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_138_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_1353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_51_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_224_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09259_ _04054_ _04360_ _04378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_182_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_33_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12270_ _01298_ clknet_leaf_232_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[31\]\[23\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_182_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11221_ _00287_ clknet_leaf_81_wb_clk_i soc.video_generator_1.h_count\[2\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_175_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_218_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_136_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6100 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11152_ _00218_ clknet_leaf_166_wb_clk_i soc.ram_encoder_0.output_bits_left\[4\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_175_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6111 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_136_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6122 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6133 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_175_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10103_ soc.ram_encoder_0.request_data_out\[5\] _04930_ _04953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_1_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6144 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6155 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_7_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11083_ _00149_ clknet_leaf_283_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[13\]\[21\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_6166 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_5432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6177 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_191_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10034_ soc.ram_encoder_0.request_address\[3\] soc.ram_encoder_0.address\[3\] _04900_
+ _04903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_6199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_1384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4720 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_208_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4731 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_114_1357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4742 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4753 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4764 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4775 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4786 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4797 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_229_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11985_ _01044_ clknet_leaf_144_wb_clk_i soc.ram_data_out\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_17_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10936_ soc.spi_video_ram_1.write_fifo.fifo_mem\[8\]\[24\] _04067_ _05430_ _05457_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_90_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_231_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_220_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10867_ _01713_ _05222_ _05412_ _05420_ _01340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_13_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_31_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_203_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10798_ _05383_ _01308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_173_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11419_ _00485_ clknet_leaf_187_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[30\]\[0\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_99_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_193_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_173_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_140_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06960_ _02609_ _02611_ _02616_ _02619_ _02620_ _02621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_67_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_214_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05911_ _01670_ soc.cpu.ALU.x\[13\] _01806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_95_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06891_ _02555_ _02556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_227_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08630_ _02157_ soc.spi_video_ram_1.write_fifo.fifo_mem\[30\]\[18\] _04011_ _04020_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_05842_ _01618_ soc.cpu.AReg.data\[9\] _01718_ soc.ram_data_out\[9\] _01741_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_23_1752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_243_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08561_ _03983_ _00470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_130_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_214_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05773_ _01561_ _01675_ _01676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_70_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xclkbuf_leaf_183_wb_clk_i clknet_5_29_0_wb_clk_i clknet_leaf_183_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_07512_ soc.spi_video_ram_1.write_fifo.fifo_mem\[29\]\[26\] _03160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_165_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08492_ _02143_ soc.spi_video_ram_1.write_fifo.fifo_mem\[28\]\[11\] _03945_ _03947_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_74_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_208_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_243_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_112_wb_clk_i clknet_opt_4_0_wb_clk_i clknet_leaf_112_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_07443_ _03088_ _03089_ _03090_ _03091_ _02929_ _03092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_165_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_210_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_206_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_221_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07374_ _02971_ soc.spi_video_ram_1.write_fifo.fifo_mem\[16\]\[11\] _03023_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_143_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09113_ _02173_ soc.spi_video_ram_1.write_fifo.fifo_mem\[20\]\[26\] _04258_ _04287_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06325_ _02178_ _00040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_198_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09044_ _01379_ _04248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_11_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06256_ soc.spi_video_ram_1.fifo_in_data\[6\] _02132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_135_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_190_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06187_ _01463_ _01516_ _02074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_219_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_191_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09946_ soc.ram_encoder_0.toggled_sram_sck _04834_ _04847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_89_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4005 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4016 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09877_ soc.rom_encoder_0.request_data_out\[14\] _04742_ _04794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_4027 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4038 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4049 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08828_ _02157_ soc.spi_video_ram_1.write_fifo.fifo_mem\[23\]\[18\] _04109_ _04131_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_3315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_246_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_230_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08759_ _04093_ _00558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_233_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_73_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1902 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1913 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11770_ _00831_ clknet_leaf_89_wb_clk_i soc.spi_video_ram_1.read_value\[0\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_246_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_198_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1924 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_213_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1946 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_202_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1957 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10721_ _05341_ _01273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1968 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1979 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_186_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10652_ _05304_ _01241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_41_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_221_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_186_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10583_ net80 _05261_ _05201_ _05265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_155_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_142_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12322_ _01350_ clknet_leaf_222_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[8\]\[1\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_196_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12253_ _01281_ clknet_leaf_210_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[31\]\[6\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_177_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_1413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11204_ _00270_ clknet_leaf_5_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[11\]\[14\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_107_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_190_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_12184_ _01212_ net87 net80 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_123_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11135_ _00201_ clknet_leaf_8_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[14\]\[15\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_68_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_237_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11066_ _00132_ clknet_leaf_260_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[13\]\[4\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_5251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_23_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_209_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10017_ soc.ram_encoder_0.request_data_out\[11\] soc.ram_encoder_0.data_out\[11\]
+ _04889_ _04894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_5284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_5295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_110_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_225_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_188_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_149_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_4583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_149_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3860 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3871 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3882 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3893 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11968_ _01027_ clknet_leaf_183_wb_clk_i soc.ram_encoder_0.request_address\[5\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_91_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10919_ _05448_ _01364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_225_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11899_ _00958_ clknet_leaf_234_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[3\]\[25\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_20_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_207_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_9_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_199_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06110_ _01921_ _02002_ _02003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_07090_ _02739_ _02743_ _02589_ _02746_ _02747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_67_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06041_ _01932_ _01933_ _01934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_246_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_86_1532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09800_ _02111_ _02456_ _02450_ _04732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_114_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07992_ soc.spi_video_ram_1.write_fifo.fifo_mem\[28\]\[18\] soc.spi_video_ram_1.write_fifo.fifo_mem\[29\]\[18\]
+ soc.spi_video_ram_1.write_fifo.fifo_mem\[30\]\[18\] soc.spi_video_ram_1.write_fifo.fifo_mem\[31\]\[18\]
+ _02717_ _02714_ _03632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_214_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09731_ soc.ram_encoder_0.output_buffer\[19\] _03814_ _03788_ soc.ram_encoder_0.request_data_out\[15\]
+ _03817_ _04693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_132_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06943_ _02580_ _02587_ _02595_ _02603_ _02604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_80_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09662_ _04641_ _00914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06874_ _01380_ _02540_ _02519_ _02543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_132_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08613_ _03998_ _04011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_05825_ _01693_ _01723_ _01725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09593_ soc.rom_encoder_0.input_buffer\[1\] _04586_ _04553_ _04597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_215_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08544_ _03974_ _00462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_242_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05756_ _01561_ _01659_ _01660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_54_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08475_ _02126_ soc.spi_video_ram_1.write_fifo.fifo_mem\[28\]\[3\] _03934_ _03938_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_05687_ _01593_ _01594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_24_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_211_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07426_ soc.spi_video_ram_1.write_fifo.fifo_mem\[0\]\[27\] soc.spi_video_ram_1.write_fifo.fifo_mem\[1\]\[27\]
+ soc.spi_video_ram_1.write_fifo.fifo_mem\[2\]\[27\] soc.spi_video_ram_1.write_fifo.fifo_mem\[3\]\[27\]
+ _03054_ _02690_ _03075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_11_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07357_ _02573_ soc.spi_video_ram_1.write_fifo.fifo_mem\[29\]\[28\] _03007_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_13_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06308_ soc.spi_video_ram_1.fifo_in_address\[7\] _02167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_109_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xcaravel_hack_soc_106 io_oeb[28] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_164_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07288_ soc.spi_video_ram_1.write_fifo.fifo_mem\[0\]\[10\] soc.spi_video_ram_1.write_fifo.fifo_mem\[1\]\[10\]
+ soc.spi_video_ram_1.write_fifo.fifo_mem\[2\]\[10\] soc.spi_video_ram_1.write_fifo.fifo_mem\[3\]\[10\]
+ _02893_ _02895_ _02938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_104_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xcaravel_hack_soc_117 io_out[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xcaravel_hack_soc_128 la_data_out[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xclkbuf_leaf_80_wb_clk_i clknet_5_10_0_wb_clk_i clknet_leaf_80_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
Xcaravel_hack_soc_139 la_data_out[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_178_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09027_ _03434_ _04224_ _04237_ _00682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_191_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06239_ _02113_ soc.spi_video_ram_1.write_fifo.fifo_mem\[18\]\[0\] _02120_ _02121_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_145_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_191_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_46_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_219_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09929_ soc.ram_encoder_0.toggled_sram_sck _04832_ _04833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_172_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_213_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3101 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3112 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_207_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3123 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3134 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_171_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3145 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_65_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3156 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3167 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3178 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11822_ _00881_ clknet_leaf_32_wb_clk_i soc.spi_video_ram_1.write_fifo.read_pointer\[4\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1710 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_199_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1721 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1732 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1743 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11753_ _00814_ clknet_leaf_295_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[4\]\[26\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1765 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1776 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1787 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10704_ _02256_ soc.spi_video_ram_1.write_fifo.fifo_mem\[29\]\[19\] _05321_ _05333_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_42_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1798 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11684_ _00745_ clknet_leaf_143_wb_clk_i soc.spi_video_ram_1.fifo_in_data\[2\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_201_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_1491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_204_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10635_ soc.spi_video_ram_1.write_fifo.fifo_mem\[19\]\[16\] soc.spi_video_ram_1.fifo_in_address\[0\]
+ _05289_ _05296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_126_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_220_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10566_ net90 soc.hack_clk_strobe _05254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_154_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12305_ _01333_ clknet_leaf_148_wb_clk_i soc.ram_encoder_0.data_out\[0\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_115_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10497_ _05172_ _05210_ _05211_ _01178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_170_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_12236_ _01264_ clknet_leaf_72_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[29\]\[18\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_108_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_123_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12167_ _01195_ clknet_leaf_168_wb_clk_i soc.ram_encoder_0.address\[12\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_2_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_150_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_155_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11118_ _00184_ clknet_leaf_43_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[12\]\[27\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_231_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12098_ _01126_ net86 soc.cpu.ALU.x\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_81_1484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_211_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_5070 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11049_ _00115_ clknet_leaf_77_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[0\]\[16\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_77_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5081 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xinput7 io_in[18] net7 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XTAP_5092 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_49_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05610_ _01469_ _01518_ _01519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_224_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06590_ _02338_ _00145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_229_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_244_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05541_ _01406_ _01443_ _01448_ _01450_ _01451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_162_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08260_ _02500_ _03777_ _03817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_60_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05472_ soc.spi_video_ram_1.state_sram_clk_counter\[7\] soc.spi_video_ram_1.state_sram_clk_counter\[6\]
+ soc.spi_video_ram_1.state_sram_clk_counter\[5\] soc.spi_video_ram_1.state_sram_clk_counter\[4\]
+ _01388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_123_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07211_ soc.spi_video_ram_1.write_fifo.fifo_mem\[12\]\[8\] soc.spi_video_ram_1.write_fifo.fifo_mem\[13\]\[8\]
+ soc.spi_video_ram_1.write_fifo.fifo_mem\[14\]\[8\] soc.spi_video_ram_1.write_fifo.fifo_mem\[15\]\[8\]
+ _02575_ _02578_ _02863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_144_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_193_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_53_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08191_ _03761_ _00322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_105_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07142_ soc.spi_video_ram_1.write_fifo.fifo_mem\[24\]\[4\] soc.spi_video_ram_1.write_fifo.fifo_mem\[25\]\[4\]
+ soc.spi_video_ram_1.write_fifo.fifo_mem\[26\]\[4\] soc.spi_video_ram_1.write_fifo.fifo_mem\[27\]\[4\]
+ _02769_ _02770_ _02798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_203_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_173_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07073_ _02716_ _02721_ _02731_ _02568_ _02732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_195_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_156_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06024_ _01844_ _01846_ _01917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_126_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_236_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_177_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07975_ _03606_ _03615_ _03616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_60_1524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_228_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09714_ _02480_ _02481_ _02485_ _04679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_5_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06926_ _02583_ _02584_ _02586_ _02587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_210_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06857_ _02526_ _02527_ _00223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09645_ soc.rom_encoder_0.data_out\[10\] soc.rom_encoder_0.request_data_out\[10\]
+ _04621_ _04631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_83_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05808_ _01705_ _01708_ _01709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_76_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09576_ _04584_ _04585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_243_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06788_ soc.rom_encoder_0.output_buffer\[17\] _02455_ _02461_ _02466_ _02467_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XTAP_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_184_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08527_ _03964_ _00455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05739_ _01640_ _01573_ _01643_ _01644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_19_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_2_0_0_wb_clk_i clknet_0_wb_clk_i clknet_2_0_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_208_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08458_ soc.spi_video_ram_1.fifo_in_address\[10\] _03927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_180_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07409_ _02941_ soc.spi_video_ram_1.write_fifo.fifo_mem\[7\]\[11\] _03058_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_08389_ _03890_ _00391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_221_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10420_ _02270_ soc.spi_video_ram_1.write_fifo.fifo_mem\[6\]\[26\] _05123_ _05152_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_87_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10351_ _01752_ _05103_ _05115_ _01129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_152_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_30_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10282_ soc.rom_loader.current_address\[0\] _01119_ _05072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_105_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12021_ _01080_ clknet_leaf_246_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[5\]\[9\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_105_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_219_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_286_wb_clk_i clknet_5_5_0_wb_clk_i clknet_leaf_286_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_234_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_215_wb_clk_i clknet_5_21_0_wb_clk_i clknet_leaf_215_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_66_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_246_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_234_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_206_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11805_ _00865_ clknet_leaf_295_wb_clk_i soc.spi_video_ram_1.fifo_in_address\[8\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_226_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_230_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_11736_ _00797_ clknet_leaf_246_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[4\]\[9\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_14_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_186_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11667_ _00728_ clknet_leaf_66_wb_clk_i soc.spi_video_ram_1.state_counter\[6\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_70_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10618_ soc.spi_video_ram_1.write_fifo.fifo_mem\[19\]\[8\] _02407_ _05278_ _05287_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_11598_ _00664_ clknet_leaf_212_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[21\]\[5\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_155_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_183_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10549_ _05222_ _01199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_122_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_143_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_157_1316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_237_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12219_ _01247_ clknet_leaf_224_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[29\]\[1\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_123_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07760_ _02712_ _03404_ _03405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_38_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_237_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_211_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06711_ soc.spi_video_ram_1.write_fifo.fifo_mem\[14\]\[9\] _02409_ _02391_ _02410_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_07691_ _02893_ soc.spi_video_ram_1.write_fifo.fifo_mem\[22\]\[24\] _03336_ _02592_
+ _03337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_246_1609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09430_ _04473_ _04482_ _04483_ _00840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06642_ _02140_ soc.spi_video_ram_1.write_fifo.fifo_mem\[12\]\[10\] _02368_ _02369_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_92_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_225_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_18_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09361_ soc.spi_video_ram_1.state_sram_clk_counter\[1\] _04432_ _04435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_1679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06573_ soc.spi_video_ram_1.write_fifo.fifo_mem\[13\]\[10\] _02237_ _02328_ _02329_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xclkbuf_leaf_19_wb_clk_i clknet_5_2_0_wb_clk_i clknet_leaf_19_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_08312_ _02153_ soc.spi_video_ram_1.write_fifo.fifo_mem\[1\]\[16\] _03842_ _03849_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_90_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05524_ _01435_ _01436_ _01396_ _00009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_209_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09292_ _04396_ _00788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_107_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_220_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_12 _02110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08243_ soc.ram_encoder_0.output_buffer\[12\] _02563_ _03804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_138_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08174_ _02159_ soc.spi_video_ram_1.write_fifo.fifo_mem\[10\]\[19\] _03743_ _03753_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_146_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07125_ _02736_ _02775_ _02780_ _02602_ _02781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_192_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07056_ soc.spi_video_ram_1.write_fifo.fifo_mem\[16\]\[2\] soc.spi_video_ram_1.write_fifo.fifo_mem\[17\]\[2\]
+ soc.spi_video_ram_1.write_fifo.fifo_mem\[18\]\[2\] soc.spi_video_ram_1.write_fifo.fifo_mem\[19\]\[2\]
+ _02713_ _02714_ _02715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_134_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_192_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_6507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06007_ _01893_ _01894_ _01899_ _01900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_6518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_6529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_102_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_5806 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_216_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5817 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5828 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5839 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_102_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_229_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_214_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07958_ _02736_ _03598_ _03599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_233_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_1444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06909_ _02569_ _02570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_07889_ _02971_ soc.spi_video_ram_1.write_fifo.fifo_mem\[4\]\[21\] _03531_ _02927_
+ _03532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_99_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_216_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09628_ _04622_ _00899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_43_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09559_ _04570_ _04571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_58_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_227_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_212_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_178_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_196_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11521_ _00587_ clknet_leaf_307_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[23\]\[15\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_134_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_106_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_211_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_200_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11452_ _00518_ clknet_leaf_53_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[15\]\[4\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10403_ _05143_ _01153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_11383_ _00449_ clknet_leaf_270_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[28\]\[22\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_125_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10334_ _01613_ _05103_ _05106_ _01121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_180_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_139_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10265_ _02272_ soc.spi_video_ram_1.write_fifo.fifo_mem\[5\]\[27\] _05041_ _05061_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_133_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12004_ _01063_ clknet_leaf_164_wb_clk_i soc.ram_encoder_0.initializing_step\[4\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_191_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10196_ soc.hack_clock_0.counter\[3\] _05020_ _05023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_121_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_94_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_219_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_235_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_169_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_207_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2060 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_146_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2071 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2082 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2093 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_202_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11719_ _00780_ clknet_leaf_283_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[9\]\[21\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_148_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_187_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_238_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xinput10 io_in[23] net10 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_204_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput21 la_data_in[12] net21 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput32 la_data_in[22] net32 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput43 la_data_in[7] net43 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_122_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_174_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_196_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xclkbuf_leaf_137_wb_clk_i clknet_5_24_0_wb_clk_i clknet_leaf_137_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_116_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_131_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08930_ soc.spi_video_ram_1.write_fifo.fifo_mem\[22\]\[7\] _02405_ _04178_ _04186_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_115_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_1387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08861_ soc.spi_video_ram_1.write_fifo.fifo_mem\[25\]\[4\] _02399_ _04144_ _04149_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_112_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_233_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07812_ _02767_ _03449_ _03456_ _02719_ _03457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_08792_ _02122_ soc.spi_video_ram_1.write_fifo.fifo_mem\[23\]\[1\] _04110_ _04112_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_84_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_215_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07743_ _02712_ _03387_ _03388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_42_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07674_ soc.spi_video_ram_1.write_fifo.fifo_mem\[5\]\[14\] _03320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_203_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_168_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09413_ _02443_ _02441_ _04459_ _02460_ _02445_ _04470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_06625_ _02124_ soc.spi_video_ram_1.write_fifo.fifo_mem\[12\]\[2\] _02357_ _02360_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_12_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09344_ _02270_ soc.spi_video_ram_1.write_fifo.fifo_mem\[4\]\[26\] _04394_ _04423_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06556_ soc.spi_video_ram_1.write_fifo.fifo_mem\[13\]\[2\] _02221_ _02317_ _02320_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_240_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_221_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_178_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05507_ _01420_ soc.spi_video_ram_1.state_sram_clk_counter\[7\] soc.spi_video_ram_1.state_sram_clk_counter\[1\]
+ _01421_ _01422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_181_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09275_ _04065_ _04360_ _04386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_139_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06487_ _02122_ soc.spi_video_ram_1.write_fifo.fifo_mem\[0\]\[1\] _02279_ _02281_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_32_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_222_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08226_ soc.ram_encoder_0.output_buffer\[4\] _03781_ _03789_ soc.ram_encoder_0.request_data_out\[0\]
+ _03790_ _03791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_33_1743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_14_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_180_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08157_ _03744_ _00305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_193_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07108_ soc.spi_video_ram_1.write_fifo.fifo_mem\[28\]\[3\] soc.spi_video_ram_1.write_fifo.fifo_mem\[29\]\[3\]
+ soc.spi_video_ram_1.write_fifo.fifo_mem\[30\]\[3\] soc.spi_video_ram_1.write_fifo.fifo_mem\[31\]\[3\]
+ _02764_ _02723_ _02765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_08088_ _03703_ _00277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_162_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07039_ _02597_ soc.spi_video_ram_1.write_fifo.fifo_mem\[4\]\[2\] _02698_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_6315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10050_ soc.ram_encoder_0.request_address\[11\] soc.ram_encoder_0.address\[11\] _04879_
+ _04911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_62_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4902 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_102_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_114_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4913 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4924 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4935 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4946 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4957 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_4968 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4979 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_217_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10952_ _00018_ clknet_leaf_247_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[18\]\[6\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_113_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_244_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_186_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10883_ _02539_ _05221_ _05411_ _05428_ _01348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_147_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_189_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_199_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_197_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_11_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11504_ _00570_ clknet_leaf_293_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[24\]\[27\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_106_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_199_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11435_ _00501_ clknet_leaf_26_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[30\]\[16\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_125_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_230_wb_clk_i clknet_5_16_0_wb_clk_i clknet_leaf_230_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_67_1316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_197_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11366_ _00432_ clknet_leaf_175_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[28\]\[5\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_125_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10317_ soc.rom_loader.current_address\[12\] _05094_ _05095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_4_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_1319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11297_ _00363_ clknet_leaf_242_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[1\]\[23\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_152_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10248_ _05052_ _01089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_152_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10179_ _05003_ _05008_ _05010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_39_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_212_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_234_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06410_ _02228_ _00075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07390_ _02767_ _03033_ _03038_ _02831_ _03039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_72_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_222_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_203_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06341_ _02188_ _00046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_163_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09060_ _02213_ soc.spi_video_ram_1.write_fifo.fifo_mem\[20\]\[0\] _04259_ _04260_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_30_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_318_wb_clk_i clknet_5_0_0_wb_clk_i clknet_leaf_318_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_72_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06272_ soc.spi_video_ram_1.fifo_in_data\[11\] _02143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_176_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08011_ soc.spi_video_ram_1.write_fifo.fifo_mem\[16\]\[17\] soc.spi_video_ram_1.write_fifo.fifo_mem\[17\]\[17\]
+ soc.spi_video_ram_1.write_fifo.fifo_mem\[18\]\[17\] soc.spi_video_ram_1.write_fifo.fifo_mem\[19\]\[17\]
+ _02681_ _02758_ _03650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_162_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_1438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_200_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09962_ _04857_ _04848_ _04858_ _00997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_176_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08913_ _02388_ _04175_ _04176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09893_ net53 _04804_ _04806_ _00980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08844_ _03927_ _04110_ _04139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_230_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_135_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_131_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05987_ soc.boot_loading_offset\[3\] _01877_ _01879_ _01880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_08775_ _04101_ _00566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_61_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_34_wb_clk_i clknet_5_9_0_wb_clk_i clknet_leaf_34_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_2807 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07726_ _02703_ soc.spi_video_ram_1.write_fifo.fifo_mem\[13\]\[24\] _03371_ _02741_
+ _03372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_2818 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2829 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_226_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07657_ _02581_ _03299_ _03302_ _03303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_207_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_228_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06608_ soc.spi_video_ram_1.write_fifo.fifo_mem\[13\]\[25\] _02268_ _02316_ _02349_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_13_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07588_ _03233_ _03234_ _02976_ _03235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_90_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_185_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06539_ _02307_ _00125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09327_ _04414_ _00805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_182_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09258_ _03308_ _04375_ _04377_ _00773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_08209_ soc.ram_encoder_0.initializing_step\[0\] _02550_ _03777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_154_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09189_ _01459_ _04339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_181_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11220_ _00286_ clknet_5_10_0_wb_clk_i soc.video_generator_1.h_count\[1\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_49_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_175_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11151_ _00217_ clknet_leaf_126_wb_clk_i net67 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_6101 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_134_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6112 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6123 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10102_ _01395_ _04952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_6134 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11082_ _00148_ clknet_leaf_48_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[13\]\[20\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_6145 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6156 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6167 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6178 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10033_ _04902_ _01024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_6189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_216_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4710 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4721 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4732 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4743 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4754 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4765 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4776 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_4787 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4798 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11984_ _01043_ clknet_leaf_155_wb_clk_i soc.ram_data_out\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_40_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_245_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_216_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10935_ _05456_ _01372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_166_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_232_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_177_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10866_ soc.ram_encoder_0.data_out\[7\] _05420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_204_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_207_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_185_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_242_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10797_ _02225_ soc.spi_video_ram_1.write_fifo.fifo_mem\[7\]\[4\] _05378_ _05383_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XPHY_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_173_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_185_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11418_ _00484_ clknet_leaf_296_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[2\]\[28\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_160_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_67_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_158_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_126_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11349_ _00415_ clknet_leaf_23_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[27\]\[17\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_98_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_234_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05910_ _01786_ _01805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_06890_ _01379_ _02548_ _02554_ _02555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
XFILLER_79_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_239_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05841_ _01702_ _01739_ _01740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_12_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_55_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_236_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05772_ _01673_ _01674_ _01675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_08560_ _02149_ soc.spi_video_ram_1.write_fifo.fifo_mem\[2\]\[14\] _03978_ _03983_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_78_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_208_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07511_ _02744_ soc.spi_video_ram_1.write_fifo.fifo_mem\[30\]\[26\] _03158_ _02908_
+ _03159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_08491_ _03946_ _00437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_235_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07442_ _02926_ soc.spi_video_ram_1.write_fifo.fifo_mem\[17\]\[27\] _03024_ _03091_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_90_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_165_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_167_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_245_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_22_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07373_ _03021_ soc.spi_video_ram_1.write_fifo.fifo_mem\[19\]\[11\] _02614_ _03022_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_182_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09112_ _04286_ _00718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06324_ _02177_ soc.spi_video_ram_1.write_fifo.fifo_mem\[18\]\[28\] _02119_ _02178_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_52_1448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_152_wb_clk_i clknet_5_30_0_wb_clk_i clknet_leaf_152_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_191_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09043_ soc.spi_video_ram_1.write_fifo.read_pointer\[1\] _04246_ _04247_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__and2_1
X_06255_ _02131_ _00017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_163_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06186_ _01460_ _02072_ _02073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_150_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_176_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_46_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_104_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09945_ soc.ram_encoder_0.input_buffer\[0\] _04846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_132_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_213_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_246_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09876_ _04787_ _04793_ _00976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_150_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4006 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4017 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4028 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4039 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08827_ _04130_ _00589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08758_ soc.spi_video_ram_1.write_fifo.fifo_mem\[24\]\[15\] _04054_ _04087_ _04093_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_2615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_241_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_227_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07709_ _02679_ _03354_ _03355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_2_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1903 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1914 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08689_ _03312_ _04046_ _04053_ _00528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_53_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1925 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1936 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1947 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10720_ _02272_ soc.spi_video_ram_1.write_fifo.fifo_mem\[29\]\[27\] _05321_ _05341_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_81_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_214_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_159_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1958 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1969 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_126_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_161_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10651_ soc.spi_video_ram_1.write_fifo.fifo_mem\[19\]\[24\] _04067_ _05277_ _05304_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_142_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_224_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10582_ _01632_ _05261_ _05264_ _01211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_210_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_167_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12321_ _01349_ clknet_leaf_191_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[8\]\[0\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_126_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_214_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_177_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_182_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_237_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12252_ _01280_ clknet_leaf_178_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[31\]\[5\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_218_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_159_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11203_ _00269_ clknet_leaf_12_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[11\]\[13\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12183_ _01211_ net87 net79 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_237_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11134_ _00200_ clknet_leaf_310_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[14\]\[14\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_1_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_235_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11065_ _00131_ clknet_leaf_262_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[13\]\[3\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_114_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_5230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10016_ _04893_ _01016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_81_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_218_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3850 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_151_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3861 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3872 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_1404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_217_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3883 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3894 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11967_ _01026_ clknet_leaf_147_wb_clk_i soc.ram_encoder_0.request_address\[4\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_17_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_220_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10918_ soc.spi_video_ram_1.write_fifo.fifo_mem\[8\]\[15\] _04054_ _05442_ _05448_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_233_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11898_ _00957_ clknet_leaf_298_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[3\]\[24\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_149_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10849_ _05410_ _01332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_203_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_200_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_145_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06040_ soc.video_generator_1.v_count\[4\] _01897_ _01852_ _01933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_12_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xclkbuf_3_2_0_wb_clk_i clknet_2_1_0_wb_clk_i clknet_3_2_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_5_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07991_ _02678_ _03630_ _03631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_114_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09730_ _04677_ _04691_ _04692_ _01381_ _00931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_06942_ _02596_ _02599_ _02602_ _02603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_132_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_45_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_227_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09661_ _04640_ soc.rom_encoder_0.request_address\[0\] _04632_ _04641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_28_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_214_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06873_ _02541_ _02542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_94_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_243_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08612_ _04010_ _00494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05824_ _01662_ _01691_ _01723_ _01724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_09592_ soc.rom_encoder_0.input_buffer\[5\] _04596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_83_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_209_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05755_ _01657_ _01658_ _01659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_08543_ _02132_ soc.spi_video_ram_1.write_fifo.fifo_mem\[2\]\[6\] _03967_ _03974_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_82_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_208_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_243_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_211_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05686_ soc.cpu.instruction\[15\] soc.cpu.instruction\[5\] _01593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_39_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08474_ _03937_ _00429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_93_1559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_196_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_210_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07425_ _02831_ _03073_ _03074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_165_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_23_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07356_ _02903_ soc.spi_video_ram_1.write_fifo.fifo_mem\[30\]\[28\] _02646_ _03006_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_109_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_52_1278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06307_ _02166_ _00034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_108_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07287_ _02831_ _02930_ _02936_ _02937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
Xcaravel_hack_soc_107 io_oeb[29] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_40_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xcaravel_hack_soc_118 io_out[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xcaravel_hack_soc_129 la_data_out[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_09026_ _04065_ _04225_ _04237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06238_ _02119_ _02120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_156_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_219_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_145_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06169_ _01994_ soc.spi_video_ram_1.read_value\[0\] _02062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_6_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_65_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09928_ soc.ram_encoder_0.request_write _02503_ _04831_ _04832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_150_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09859_ _04752_ _04780_ _00972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_8_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3102 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3113 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3124 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3135 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3146 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_233_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3157 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3168 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11821_ _00880_ clknet_leaf_32_wb_clk_i soc.spi_video_ram_1.write_fifo.read_pointer\[3\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3179 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1700 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_164_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1711 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1722 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1733 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_202_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11752_ _00813_ clknet_leaf_287_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[4\]\[25\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_14_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1744 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_215_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1755 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_18_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1766 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_186_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10703_ _05332_ _01264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1788 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_183_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11683_ _00744_ clknet_leaf_145_wb_clk_i soc.spi_video_ram_1.fifo_in_data\[1\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_14_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1799 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10634_ _05295_ _01232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_122_1413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_204_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_1446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10565_ _03714_ _05253_ _01205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_10_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_196_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12304_ _01332_ clknet_leaf_274_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[7\]\[28\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10496_ soc.cpu.PC.in\[12\] _05188_ _05201_ _05211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_120_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_12235_ _01263_ clknet_leaf_73_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[29\]\[17\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_108_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_190_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_233_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12166_ _01194_ clknet_leaf_153_wb_clk_i soc.ram_encoder_0.address\[11\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_155_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11117_ _00183_ clknet_leaf_279_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[12\]\[26\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_110_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_12097_ _01125_ net86 soc.cpu.ALU.x\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_211_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_209_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5060 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_133_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11048_ _00114_ clknet_leaf_321_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[0\]\[15\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_5071 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xinput8 io_in[19] net8 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_188_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_5082 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_225_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5093 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_209_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05540_ _01407_ _01449_ _01450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_75_1245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_221_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_178_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2990 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05471_ soc.spi_video_ram_1.state_sram_clk_counter\[8\] _01387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_162_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_18_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07210_ _02583_ _02861_ _02862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_08190_ _02175_ soc.spi_video_ram_1.write_fifo.fifo_mem\[10\]\[27\] _03731_ _03761_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_07141_ _02571_ _02796_ _02586_ _02797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_105_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_238_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07072_ _02583_ _02724_ _02730_ _02586_ _02731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_118_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_220_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06023_ _01908_ _01914_ _01915_ _01916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_133_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_1314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_160_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07974_ _03608_ _03610_ _03612_ _03614_ _02568_ _03615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_5_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09713_ _02549_ _02553_ _04677_ _04678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_45_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06925_ _02585_ _02586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_132_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_132_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09644_ _04630_ _00907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_67_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06856_ soc.rom_encoder_0.output_bits_left\[2\] _02513_ _02527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_56_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_228_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_215_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_186_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_1749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05807_ _01706_ _01707_ _01708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_110_1350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09575_ soc.rom_encoder_0.toggled_sram_sck _04566_ _04584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_83_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06787_ _02443_ _02465_ _02466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_167_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08526_ _02177_ soc.spi_video_ram_1.write_fifo.fifo_mem\[28\]\[28\] _03933_ _03964_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_05738_ net80 _01642_ _01575_ soc.gpio_i_stored\[3\] _01573_ _01643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_54_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_211_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_168_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08457_ _03926_ _00423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05669_ soc.cpu.AReg.data\[1\] _01566_ _01577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_36_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07408_ _02941_ soc.spi_video_ram_1.write_fifo.fifo_mem\[5\]\[11\] _03056_ _03057_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_184_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08388_ soc.spi_video_ram_1.write_fifo.fifo_mem\[26\]\[22\] _02262_ _03865_ _03890_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_17_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_137_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07339_ _02712_ soc.spi_video_ram_1.write_fifo.fifo_mem\[4\]\[28\] _02741_ _02989_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_109_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10350_ soc.cpu.ALU.x\[9\] _05109_ _05115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_191_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09009_ _03291_ _04224_ _04228_ _00673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_10281_ _05070_ _05071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_139_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_69_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_191_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12020_ _01079_ clknet_leaf_228_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[5\]\[8\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_133_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_215_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_238_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_19_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_207_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_189_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xclkbuf_leaf_255_wb_clk_i clknet_5_18_0_wb_clk_i clknet_leaf_255_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_46_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_98_1278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_185_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11804_ _00864_ clknet_leaf_286_wb_clk_i soc.spi_video_ram_1.fifo_in_address\[7\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_203_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_187_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11735_ _00796_ clknet_leaf_228_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[4\]\[8\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_163_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_204_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_187_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11666_ _00727_ clknet_leaf_83_wb_clk_i soc.spi_video_ram_1.state_counter\[5\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_126_1390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_50_1749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10617_ _05286_ _01224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_11597_ _00663_ clknet_leaf_132_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[21\]\[4\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_183_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_239_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10548_ _05224_ _01198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_115_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_170_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10479_ soc.cpu.PC.in\[8\] _05188_ _05173_ _05198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_29_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12218_ _01246_ clknet_leaf_187_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[29\]\[0\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_48_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_123_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_170_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_151_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12149_ _01177_ net88 soc.cpu.PC.REG.data\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_42_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06710_ soc.spi_video_ram_1.fifo_in_data\[9\] _02409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_07690_ _02612_ _03335_ _03336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_53_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_25_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06641_ _02355_ _02368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_168_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_129_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09360_ _04432_ _04434_ _00818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_244_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_240_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06572_ _02315_ _02328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_166_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_5_23_0_wb_clk_i clknet_4_11_0_wb_clk_i clknet_5_23_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_181_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08311_ _03848_ _00355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_75_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_05523_ soc.spi_video_ram_1.initialized soc.spi_video_ram_1.start_read soc.spi_video_ram_1.current_state\[2\]
+ _01408_ _01436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_21_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09291_ _02213_ soc.spi_video_ram_1.write_fifo.fifo_mem\[4\]\[0\] _04395_ _04396_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_61_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_13 soc.cpu.AReg.data\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_166_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08242_ soc.ram_encoder_0.output_buffer\[8\] _03781_ _03789_ soc.ram_encoder_0.request_data_out\[4\]
+ _03802_ _03803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_53_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_59_wb_clk_i clknet_5_13_0_wb_clk_i clknet_leaf_59_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_08173_ _03752_ _00313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_203_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07124_ _02776_ _02777_ _02589_ _02779_ _02780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_174_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_146_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07055_ _02598_ _02714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
X_06006_ _01895_ _01896_ _01898_ _01899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_66_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_161_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5807 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5818 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_114_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5829 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_130_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07957_ soc.spi_video_ram_1.write_fifo.fifo_mem\[8\]\[19\] soc.spi_video_ram_1.write_fifo.fifo_mem\[9\]\[19\]
+ soc.spi_video_ram_1.write_fifo.fifo_mem\[10\]\[19\] soc.spi_video_ram_1.write_fifo.fifo_mem\[11\]\[19\]
+ _02713_ _02737_ _03598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_87_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_116_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_210_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_244_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06908_ _00002_ _02569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_07888_ _02688_ _03530_ _03531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_28_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09627_ soc.rom_encoder_0.data_out\[1\] soc.rom_encoder_0.request_data_out\[1\] _04621_
+ _04622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06839_ _02511_ _02512_ _00220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_71_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_243_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09558_ soc.rom_encoder_0.input_bits_left\[4\] _04569_ _04570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_19_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08509_ _03955_ _00446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_24_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09489_ _01428_ _02091_ _04529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_93_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11520_ _00586_ clknet_leaf_3_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[23\]\[14\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_221_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11451_ _00517_ clknet_leaf_53_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[15\]\[3\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_201_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_137_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_165_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10402_ _02252_ soc.spi_video_ram_1.write_fifo.fifo_mem\[6\]\[17\] _05135_ _05143_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_137_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11382_ _00448_ clknet_leaf_291_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[28\]\[21\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_194_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10333_ soc.cpu.ALU.x\[1\] _05104_ _05106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_178_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_219_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10264_ _03178_ _05044_ _05060_ _01097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_65_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_234_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12003_ _01062_ clknet_leaf_163_wb_clk_i soc.ram_encoder_0.initializing_step\[3\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_156_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10195_ soc.hack_clock_0.counter\[3\] _05020_ _05022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_87_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_239_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_43_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_234_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_185_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2050 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_222_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2061 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_50_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_62_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2072 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2083 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_226_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_167_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2094 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11718_ _00779_ clknet_leaf_53_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[9\]\[20\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_30_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput11 io_in[24] net11 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_11649_ _00710_ clknet_leaf_27_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[20\]\[17\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xinput22 la_data_in[13] net22 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_128_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput33 la_data_in[23] net33 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_200_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput44 la_data_in[8] net44 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_7_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_48_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_177_wb_clk_i clknet_5_23_0_wb_clk_i clknet_leaf_177_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_08860_ _04148_ _00604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_111_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07811_ _02582_ _03452_ _03455_ _03456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_97_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_229_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_106_wb_clk_i clknet_5_14_0_wb_clk_i clknet_leaf_106_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_170_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08791_ _04111_ _00572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_85_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_226_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_211_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07742_ soc.spi_video_ram_1.write_fifo.fifo_mem\[21\]\[15\] _03387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_113_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07673_ soc.spi_video_ram_1.write_fifo.fifo_mem\[0\]\[14\] soc.spi_video_ram_1.write_fifo.fifo_mem\[1\]\[14\]
+ soc.spi_video_ram_1.write_fifo.fifo_mem\[2\]\[14\] soc.spi_video_ram_1.write_fifo.fifo_mem\[3\]\[14\]
+ _02902_ _02894_ _03319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_38_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_225_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09412_ _04468_ _02441_ _02515_ _02454_ _04469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_129_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_92_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06624_ _02359_ _00158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_20_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_241_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_179_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09343_ _04422_ _00813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_90_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06555_ _02319_ _00129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_209_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_224_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05506_ soc.spi_video_ram_1.state_sram_clk_counter\[3\] _01415_ soc.spi_video_ram_1.state_sram_clk_counter\[0\]
+ _01421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_146_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09274_ _03517_ _04375_ _04385_ _00781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_240_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06486_ _02280_ _00099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_33_1722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_194_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08225_ soc.ram_encoder_0.request_address\[7\] _02506_ _03790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_21_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08156_ _02140_ soc.spi_video_ram_1.write_fifo.fifo_mem\[10\]\[10\] _03743_ _03744_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_147_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_140_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07107_ _02763_ _02764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_134_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08087_ soc.spi_video_ram_1.write_fifo.fifo_mem\[11\]\[21\] _02260_ _03679_ _03703_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_106_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_136_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_164_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07038_ _02696_ _02697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_6305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_134_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_216_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_88_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_88_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4903 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4914 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_130_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_180_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08989_ soc.spi_video_ram_1.write_fifo.fifo_mem\[21\]\[6\] _02403_ _04210_ _04217_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_4925 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4936 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4947 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4958 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_151_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4969 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_216_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_186_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10951_ _00017_ clknet_leaf_215_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[18\]\[5\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_90_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_204_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10882_ soc.ram_encoder_0.data_out\[15\] _05428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_227_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_231_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_244_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_164_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_196_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_200_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11503_ _00569_ clknet_leaf_292_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[24\]\[26\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_157_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11434_ _00500_ clknet_leaf_309_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[30\]\[15\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_201_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11365_ _00431_ clknet_leaf_195_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[28\]\[4\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_153_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_4_wb_clk_i clknet_5_2_0_wb_clk_i clknet_leaf_4_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_99_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10316_ _05070_ _05093_ _05094_ _01114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_154_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11296_ _00362_ clknet_leaf_251_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[1\]\[22\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_140_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_191_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_270_wb_clk_i clknet_5_6_0_wb_clk_i clknet_leaf_270_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_10247_ _02254_ soc.spi_video_ram_1.write_fifo.fifo_mem\[5\]\[18\] _05041_ _05052_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_80_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10178_ _05007_ _05005_ _05009_ _03714_ _01062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_117_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_208_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_235_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_207_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_39_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_223_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_143_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_50_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_124_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06340_ _02130_ soc.spi_video_ram_1.write_fifo.fifo_mem\[17\]\[5\] _02182_ _02188_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_206_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_241_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_187_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06271_ _02142_ _00022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_72_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_204_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08010_ _03577_ _03648_ _03579_ _03649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_106_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_159_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_156_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_184_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_1406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_1488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_239_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09961_ soc.ram_encoder_0.input_buffer\[0\] _04849_ _04248_ _04858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_104_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08912_ _02116_ _04107_ _04175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_217_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_174_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09892_ _01395_ _04805_ _04806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_170_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08843_ _03237_ _04124_ _04138_ _00597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_100_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_246_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_170_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_170_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_230_1753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08774_ soc.spi_video_ram_1.write_fifo.fifo_mem\[24\]\[23\] _04065_ _04075_ _04101_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_05986_ _01869_ _01873_ _01878_ _01879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_2_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07725_ _02573_ soc.spi_video_ram_1.write_fifo.fifo_mem\[12\]\[24\] _03371_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_72_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2808 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2819 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07656_ _02574_ soc.spi_video_ram_1.write_fifo.fifo_mem\[28\]\[14\] _03301_ _02741_
+ _03302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_20_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_246_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06607_ _02348_ _00152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xclkbuf_leaf_74_wb_clk_i clknet_5_9_0_wb_clk_i clknet_leaf_74_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_213_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07587_ _02926_ soc.spi_video_ram_1.write_fifo.fifo_mem\[16\]\[25\] _03234_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_107_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_240_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09326_ _02252_ soc.spi_video_ram_1.write_fifo.fifo_mem\[4\]\[17\] _04406_ _04414_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_178_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_146_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06538_ _02173_ soc.spi_video_ram_1.write_fifo.fifo_mem\[0\]\[26\] _02278_ _02307_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_09257_ _04052_ _04375_ _04377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06469_ soc.spi_video_ram_1.fifo_in_address\[9\] _02268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_167_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_239_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08208_ _01381_ _03776_ _00324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09188_ _01589_ _04338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_193_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08139_ _02124_ soc.spi_video_ram_1.write_fifo.fifo_mem\[10\]\[2\] _03732_ _03735_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_159_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_190_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_194_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11150_ _00216_ clknet_leaf_125_wb_clk_i net66 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_6102 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6113 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10101_ _04787_ _04951_ _01042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_150_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6124 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_136_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6135 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11081_ _00147_ clknet_leaf_35_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[13\]\[19\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_6146 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6157 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_6168 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10032_ soc.ram_encoder_0.request_address\[2\] soc.ram_encoder_0.address\[2\] _04900_
+ _04902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6179 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_23_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_194_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_4700 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_114_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4711 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_49_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4722 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4733 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4744 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4755 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4766 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_217_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4777 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4788 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11983_ _01042_ clknet_leaf_158_wb_clk_i soc.ram_data_out\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_91_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4799 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_244_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_56_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xclkbuf_4_4_0_wb_clk_i clknet_3_2_0_wb_clk_i clknet_4_4_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_10934_ soc.spi_video_ram_1.write_fifo.fifo_mem\[8\]\[23\] _04065_ _05430_ _05456_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_205_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_186_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_182_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10865_ _01699_ _05222_ _05412_ _05419_ _01339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_31_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_125_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_197_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10796_ _05382_ _01307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_223_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_205_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11417_ _00483_ clknet_leaf_42_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[2\]\[27\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_197_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11348_ _00414_ clknet_leaf_19_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[27\]\[16\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_113_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_154_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11279_ _00345_ clknet_leaf_215_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[1\]\[5\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_140_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_95_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_66_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05840_ _01670_ soc.cpu.ALU.x\[9\] _01739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_212_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5990 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05771_ _01598_ soc.cpu.AReg.data\[5\] _01606_ _01674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07510_ _02903_ _03157_ _03158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_81_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08490_ _02140_ soc.spi_video_ram_1.write_fifo.fifo_mem\[28\]\[10\] _03945_ _03946_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_1_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07441_ _02752_ soc.spi_video_ram_1.write_fifo.fifo_mem\[16\]\[27\] _03090_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_222_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07372_ _02695_ _03021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_91_1465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09111_ _02171_ soc.spi_video_ram_1.write_fifo.fifo_mem\[20\]\[25\] _04258_ _04286_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_31_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06323_ soc.spi_video_ram_1.fifo_in_address\[12\] _02177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_104_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09042_ _04243_ _04245_ _04246_ _00688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_15_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06254_ _02130_ soc.spi_video_ram_1.write_fifo.fifo_mem\[18\]\[5\] _02120_ _02131_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_191_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_191_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_192_wb_clk_i clknet_5_28_0_wb_clk_i clknet_leaf_192_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_198_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06185_ _01469_ _01470_ _01463_ _02072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_209_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_176_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_172_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_121_wb_clk_i clknet_5_15_0_wb_clk_i clknet_leaf_121_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_144_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_176_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09944_ _04842_ _04844_ _04845_ _00992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_172_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09875_ soc.cpu.instruction\[13\] _04741_ _04792_ _04793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4007 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4018 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4029 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08826_ _02155_ soc.spi_video_ram_1.write_fifo.fifo_mem\[23\]\[17\] _04109_ _04130_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_6_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_3317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08757_ _04092_ _00557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05969_ soc.video_generator_1.v_count\[1\] _01862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XTAP_2605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_226_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07708_ soc.spi_video_ram_1.write_fifo.fifo_mem\[7\]\[24\] _03354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_38_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1904 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08688_ _04052_ _04048_ _04053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_187_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_242_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1926 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07639_ _02931_ soc.spi_video_ram_1.write_fifo.fifo_mem\[17\]\[14\] _03285_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1948 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1959 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_241_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10650_ _05303_ _01240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_198_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09309_ _02235_ soc.spi_video_ram_1.write_fifo.fifo_mem\[4\]\[9\] _04395_ _04405_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_10581_ net79 _05261_ _05201_ _05264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_155_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_142_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12320_ _01348_ clknet_leaf_117_wb_clk_i soc.ram_encoder_0.data_out\[15\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_161_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_202_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12251_ _01279_ clknet_leaf_140_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[31\]\[4\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_207_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11202_ _00268_ clknet_leaf_2_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[11\]\[12\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_68_1445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12182_ _01210_ net87 net78 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_123_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_1426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11133_ _00199_ clknet_leaf_11_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[14\]\[13\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_150_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11064_ _00130_ clknet_leaf_137_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[13\]\[2\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_122_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10015_ soc.ram_encoder_0.request_data_out\[10\] soc.ram_encoder_0.data_out\[10\]
+ _04889_ _04893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_5264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_149_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3840 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3851 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3862 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3873 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11966_ _01025_ clknet_leaf_146_wb_clk_i soc.ram_encoder_0.request_address\[3\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3884 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3895 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10917_ _05447_ _01363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_232_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11897_ _00956_ clknet_leaf_241_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[3\]\[23\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_92_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_204_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10848_ _02274_ soc.spi_video_ram_1.write_fifo.fifo_mem\[7\]\[28\] _05389_ _05410_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_158_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_242_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_220_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10779_ _04069_ _05359_ _05373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_121_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_220_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_158_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_195_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_1501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07990_ soc.spi_video_ram_1.write_fifo.fifo_mem\[24\]\[18\] soc.spi_video_ram_1.write_fifo.fifo_mem\[25\]\[18\]
+ soc.spi_video_ram_1.write_fifo.fifo_mem\[26\]\[18\] soc.spi_video_ram_1.write_fifo.fifo_mem\[27\]\[18\]
+ _02681_ _02758_ _03630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_218_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_101_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06941_ _02601_ _02602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_113_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_1718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09660_ soc.cpu.PC.REG.data\[0\] soc.rom_loader.current_address\[0\] _04639_ _04640_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06872_ _01379_ _02540_ _02541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_228_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08611_ _02138_ soc.spi_video_ram_1.write_fifo.fifo_mem\[30\]\[9\] _04000_ _04010_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_83_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05823_ _01689_ _01711_ _01710_ _01723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_09591_ _04594_ _04585_ _04595_ _00889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_55_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_227_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_208_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08542_ _03973_ _00461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05754_ _01598_ soc.cpu.AReg.data\[4\] _01606_ _01658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_224_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_1527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08473_ _02124_ soc.spi_video_ram_1.write_fifo.fifo_mem\[28\]\[2\] _03934_ _03937_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_05685_ _01553_ _01554_ _01555_ _01589_ _01592_ _01564_ soc.cpu.PC.in\[0\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai222_2
XFILLER_145_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07424_ _03069_ _03070_ _03071_ _03072_ _02929_ _03073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_223_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07355_ _02695_ soc.spi_video_ram_1.write_fifo.fifo_mem\[31\]\[28\] _03005_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_91_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_210_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_206_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06306_ _02165_ soc.spi_video_ram_1.write_fifo.fifo_mem\[18\]\[22\] _02119_ _02166_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xclkbuf_leaf_302_wb_clk_i clknet_5_4_0_wb_clk_i clknet_leaf_302_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_07286_ _02691_ _02933_ _02934_ _02935_ _02588_ _02936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_163_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xcaravel_hack_soc_108 io_oeb[34] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xcaravel_hack_soc_119 io_out[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_09025_ _03485_ _04224_ _04236_ _00681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_164_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06237_ _02118_ _02119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_69_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_145_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06168_ soc.spi_video_ram_1.read_value\[1\] _02061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_176_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06099_ _01970_ _01991_ _01992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_160_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_172_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09927_ soc.ram_encoder_0.current_state\[2\] _04830_ _04831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_104_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_1432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_232_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09858_ _01717_ _04740_ _04779_ _04780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3103 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3114 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08809_ _02138_ soc.spi_video_ram_1.write_fifo.fifo_mem\[23\]\[9\] _04117_ _04121_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_98_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3125 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09789_ _04724_ _00958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3136 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3147 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_185_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_227_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11820_ _00879_ clknet_leaf_47_wb_clk_i soc.spi_video_ram_1.write_fifo.read_pointer\[2\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3169 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1701 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1712 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1723 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_183_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_11751_ _00812_ clknet_leaf_302_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[4\]\[24\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_214_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_157_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1745 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1756 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_183_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1767 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10702_ _02254_ soc.spi_video_ram_1.write_fifo.fifo_mem\[29\]\[18\] _05321_ _05332_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_1778 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11682_ _00743_ clknet_leaf_186_wb_clk_i soc.spi_video_ram_1.fifo_in_data\[0\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_35_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1789 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_197_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_202_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10633_ soc.spi_video_ram_1.write_fifo.fifo_mem\[19\]\[15\] _04054_ _05289_ _05295_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_224_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10564_ soc.boot_loading_offset\[4\] _05252_ _05253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_10_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_194_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_155_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12303_ _01331_ clknet_leaf_272_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[7\]\[27\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10495_ soc.cpu.PC.REG.data\[12\] _05209_ _05210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_136_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12234_ _01262_ clknet_leaf_30_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[29\]\[16\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_108_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_151_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12165_ _01193_ clknet_leaf_151_wb_clk_i soc.ram_encoder_0.address\[10\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_151_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11116_ _00182_ clknet_leaf_286_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[12\]\[25\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_235_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_12096_ _01124_ net86 soc.cpu.ALU.x\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_150_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5050 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11047_ _00113_ clknet_leaf_321_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[0\]\[14\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_5061 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5072 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_49_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xinput9 io_in[22] net9 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XTAP_5083 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5094 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_7_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_209_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_206_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3692 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_5_13_0_wb_clk_i clknet_4_6_0_wb_clk_i clknet_5_13_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_11949_ _01008_ clknet_leaf_156_wb_clk_i soc.ram_encoder_0.request_data_out\[2\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_233_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2980 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2991 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_205_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05470_ soc.spi_video_ram_1.state_sram_clk_counter\[1\] _01386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_127_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_221_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_203_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_192_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07140_ soc.spi_video_ram_1.write_fifo.fifo_mem\[28\]\[4\] soc.spi_video_ram_1.write_fifo.fifo_mem\[29\]\[4\]
+ soc.spi_video_ram_1.write_fifo.fifo_mem\[30\]\[4\] soc.spi_video_ram_1.write_fifo.fifo_mem\[31\]\[4\]
+ _02689_ _02723_ _02796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_146_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_72_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_119_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07071_ _02725_ _02727_ _02729_ _02693_ _02707_ _02730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_06022_ _01910_ _01913_ _01915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_127_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_86_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_86_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_236_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07973_ _02571_ _03613_ _02602_ _03614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_190_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_116_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_25_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09712_ _02548_ _02554_ _04677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_151_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06924_ _00003_ _02585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_99_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_214_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09643_ soc.rom_encoder_0.data_out\[9\] soc.rom_encoder_0.request_data_out\[9\] _04621_
+ _04630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06855_ soc.rom_encoder_0.output_bits_left\[2\] _02513_ _02525_ _02526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_99_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_209_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05806_ _01598_ soc.cpu.AReg.data\[7\] _01606_ _01707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_82_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09574_ soc.rom_encoder_0.input_buffer\[0\] _04583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_43_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06786_ soc.rom_encoder_0.output_buffer\[17\] _02463_ _02464_ soc.rom_encoder_0.request_data_out\[13\]
+ _02465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_227_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_231_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_208_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08525_ _03963_ _00454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_149_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05737_ soc.cpu.AReg.data\[0\] _01572_ _01641_ _01642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_24_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_227_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_196_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08456_ soc.spi_video_ram_1.write_fifo.fifo_mem\[27\]\[25\] _02268_ _03898_ _03926_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_05668_ _01568_ _01569_ _01570_ _01571_ _01576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_23_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07407_ _02644_ soc.spi_video_ram_1.write_fifo.fifo_mem\[4\]\[11\] _03056_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_52_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08387_ _03889_ _00390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05599_ soc.spi_video_ram_1.output_buffer\[19\] _01508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_225_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_211_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07338_ _02703_ soc.spi_video_ram_1.write_fifo.fifo_mem\[5\]\[28\] _02988_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_104_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07269_ _02573_ _02919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_118_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_192_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09008_ _04052_ _04225_ _04228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_10280_ _04426_ soc.rom_loader.was_loading _05070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_164_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_156_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_120_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_76_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_8_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11803_ _00863_ clknet_leaf_265_wb_clk_i soc.spi_video_ram_1.fifo_in_address\[6\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_221_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_295_wb_clk_i clknet_5_4_0_wb_clk_i clknet_leaf_295_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_15_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_215_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_11734_ _00795_ clknet_leaf_244_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[4\]\[7\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_186_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xclkbuf_leaf_224_wb_clk_i clknet_5_23_0_wb_clk_i clknet_leaf_224_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XPHY_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_203_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11665_ _00726_ clknet_leaf_67_wb_clk_i soc.spi_video_ram_1.state_counter\[4\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_174_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10616_ soc.spi_video_ram_1.write_fifo.fifo_mem\[19\]\[7\] _02405_ _05278_ _05286_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_122_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11596_ _00662_ clknet_leaf_132_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[21\]\[3\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_127_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_204_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_196_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10547_ _05243_ _01197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_183_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10478_ soc.cpu.PC.REG.data\[8\] _05196_ _05197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_12217_ _01245_ clknet_leaf_280_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[19\]\[28\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_29_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_233_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_124_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12148_ _01176_ net88 soc.cpu.PC.REG.data\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_110_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12079_ soc.cpu.PC.in\[2\] net84 soc.cpu.AReg.data\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_111_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_133_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_238_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06640_ _02367_ _00166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_4190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_52_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_213_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_209_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06571_ _02327_ _00137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_80_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08310_ _02151_ soc.spi_video_ram_1.write_fifo.fifo_mem\[1\]\[15\] _03842_ _03848_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_127_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_55_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05522_ _01419_ _01434_ _01435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_162_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09290_ _04394_ _04395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_127_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_244_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08241_ soc.ram_encoder_0.request_address\[11\] _02505_ _03802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA_14 net25 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_193_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08172_ _02157_ soc.spi_video_ram_1.write_fifo.fifo_mem\[10\]\[18\] _03743_ _03752_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_140_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_158_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07123_ _02697_ soc.spi_video_ram_1.write_fifo.fifo_mem\[7\]\[4\] _02778_ _02723_
+ _02779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_88_1426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_99_wb_clk_i clknet_5_14_0_wb_clk_i clknet_leaf_99_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_133_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07054_ _02712_ _02713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_06005_ soc.video_generator_1.v_count\[0\] _01897_ _01898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_86_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_173_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_28_wb_clk_i clknet_5_8_0_wb_clk_i clknet_leaf_28_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_6509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_217_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_5808 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5819 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_102_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_130_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07956_ _03595_ _03596_ _03597_ _00251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_29_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06907_ _02567_ _02568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_96_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07887_ soc.spi_video_ram_1.write_fifo.fifo_mem\[5\]\[21\] _03530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_56_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_228_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_186_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06838_ soc.ram_encoder_0.output_bits_left\[2\] _02494_ _02512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09626_ _04617_ _04621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_83_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_244_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09557_ soc.rom_encoder_0.input_bits_left\[2\] _04568_ _04569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_110_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_203_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06769_ _02441_ _02446_ _02447_ _02111_ _02448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_58_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_169_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_197_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08508_ _02159_ soc.spi_video_ram_1.write_fifo.fifo_mem\[28\]\[19\] _03945_ _03955_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_180_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_184_1282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09488_ _02882_ _04528_ _00853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_223_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08439_ _03917_ _00414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_145_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_8_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_156_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_201_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_11450_ _00516_ clknet_leaf_55_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[15\]\[2\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_71_1485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10401_ _05142_ _01152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_197_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11381_ _00447_ clknet_leaf_52_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[28\]\[20\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_178_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10332_ _01589_ _05103_ _05105_ _01120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_11_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10263_ soc.spi_video_ram_1.fifo_in_address\[10\] _05045_ _05060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_2_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_3_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_12002_ _01061_ clknet_leaf_163_wb_clk_i soc.ram_encoder_0.initializing_step\[2\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_105_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10194_ _05017_ _05020_ _05021_ _01066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_238_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_228_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_34_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_210_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2040 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2051 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2062 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2073 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2084 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2095 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_99_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_245_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11717_ _00778_ clknet_leaf_32_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[9\]\[19\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_50_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11648_ _00709_ clknet_leaf_29_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[20\]\[16\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_175_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput12 io_in[25] net12 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput23 la_data_in[14] net23 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_122_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput34 la_data_in[24] net34 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput45 la_data_in[9] net45 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_122_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_239_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11579_ _00645_ clknet_leaf_276_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[22\]\[15\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_171_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_176_1749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_192_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_135_1413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07810_ _02971_ soc.spi_video_ram_1.write_fifo.fifo_mem\[4\]\[23\] _03454_ _03024_
+ _03455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_69_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_112_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_61_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08790_ _02113_ soc.spi_video_ram_1.write_fifo.fifo_mem\[23\]\[0\] _04110_ _04111_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_111_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_42_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07741_ _02704_ soc.spi_video_ram_1.write_fifo.fifo_mem\[23\]\[15\] _02958_ _03386_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_244_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_146_wb_clk_i clknet_5_28_0_wb_clk_i clknet_leaf_146_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_07672_ _02585_ _03311_ _03317_ _03318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_93_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_168_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09411_ soc.rom_encoder_0.request_address\[6\] _04468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_1423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_226_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06623_ _02122_ soc.spi_video_ram_1.write_fifo.fifo_mem\[12\]\[1\] _02357_ _02359_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_168_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_240_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09342_ _02268_ soc.spi_video_ram_1.write_fifo.fifo_mem\[4\]\[25\] _04394_ _04422_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_181_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06554_ soc.spi_video_ram_1.write_fifo.fifo_mem\[13\]\[1\] _02219_ _02317_ _02319_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_61_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05505_ _01387_ _01420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09273_ _04063_ _04360_ _04385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_90_1349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_205_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_179_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_139_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06485_ _02113_ soc.spi_video_ram_1.write_fifo.fifo_mem\[0\]\[0\] _02279_ _02280_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_08224_ _03788_ _03789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_138_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08155_ _03730_ _03743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_119_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_162_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07106_ _02644_ _02763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xclkbuf_5_6_0_wb_clk_i clknet_4_3_0_wb_clk_i clknet_5_6_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_08086_ _03702_ _00276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_134_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07037_ _02695_ _02696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_161_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_138_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4904 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4915 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08988_ _04216_ _00664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_4926 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_102_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_4937 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_180_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_4948 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_169_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07939_ soc.spi_video_ram_1.write_fifo.fifo_mem\[0\]\[20\] soc.spi_video_ram_1.write_fifo.fifo_mem\[1\]\[20\]
+ soc.spi_video_ram_1.write_fifo.fifo_mem\[2\]\[20\] soc.spi_video_ram_1.write_fifo.fifo_mem\[3\]\[20\]
+ _02764_ _02723_ _03581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_4959 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10950_ _00016_ clknet_leaf_139_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[18\]\[4\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_29_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_229_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_243_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_232_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09609_ soc.rom_encoder_0.input_buffer\[6\] _04584_ _04601_ _04608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_44_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10881_ _01834_ _05221_ _05411_ _05427_ _01347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XPHY_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_43_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_38_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_145_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_237_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_160_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_185_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_11502_ _00568_ clknet_leaf_230_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[24\]\[25\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_157_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_199_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_12_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11433_ _00499_ clknet_leaf_317_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[30\]\[14\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_240_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11364_ _00430_ clknet_leaf_138_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[28\]\[3\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_158_1435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_152_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10315_ soc.rom_loader.current_address\[11\] _05092_ _05094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_158_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_1408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_193_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11295_ _00361_ clknet_leaf_229_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[1\]\[21\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_234_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10246_ _05051_ _01088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_156_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_239_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10177_ soc.ram_encoder_0.initializing_step\[3\] _05003_ _05004_ _05008_ _05009_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_78_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_226_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_169_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_208_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_222_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06270_ _02140_ soc.spi_video_ram_1.write_fifo.fifo_mem\[18\]\[10\] _02141_ _02142_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_124_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_147_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_198_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_200_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_143_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09960_ soc.ram_encoder_0.input_buffer\[4\] _04857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_48_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08911_ _04174_ _00629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09891_ soc.rom_encoder_0.current_state\[2\] _02457_ _04614_ _04805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XTAP_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_97_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08842_ _04069_ _04110_ _04138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_44_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08773_ _04100_ _00565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_245_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_211_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05985_ _01859_ _01864_ soc.boot_loading_offset\[2\] _01878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_73_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07724_ _03139_ soc.spi_video_ram_1.write_fifo.fifo_mem\[14\]\[24\] _03369_ _02646_
+ _03370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_22_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2809 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_225_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_214_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07655_ _02902_ _03300_ _03301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_246_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_241_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_198_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06606_ soc.spi_video_ram_1.write_fifo.fifo_mem\[13\]\[24\] _02266_ _02316_ _02348_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_179_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07586_ _02920_ soc.spi_video_ram_1.write_fifo.fifo_mem\[17\]\[25\] _03233_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_25_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_209_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_80_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_224_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09325_ _04413_ _00804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06537_ _02306_ _00124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_167_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09256_ _03210_ _04375_ _04376_ _00772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_194_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06468_ _02267_ _00094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_103_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08207_ _02452_ _03771_ _03774_ _03775_ _02540_ net64 _03776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai33_1
XFILLER_21_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xclkbuf_leaf_43_wb_clk_i clknet_5_6_0_wb_clk_i clknet_leaf_43_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_194_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09187_ _01853_ _04336_ _04337_ _04317_ _00742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_06399_ soc.spi_video_ram_1.fifo_in_data\[2\] _02221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_88_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08138_ _03734_ _00296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_135_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_175_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08069_ soc.spi_video_ram_1.write_fifo.fifo_mem\[11\]\[12\] _02242_ _03691_ _03694_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_6103 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_175_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10100_ soc.ram_data_out\[4\] _04927_ _04950_ _04951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_66_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_235_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6114 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6125 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11080_ _00146_ clknet_leaf_21_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[13\]\[18\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_216_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_157_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6136 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6147 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6158 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10031_ _04901_ _01023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_6169 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_88_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_88_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4701 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_237_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4712 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_208_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4723 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_130_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4734 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_187_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4745 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4756 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4767 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4778 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4789 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11982_ _01041_ clknet_leaf_157_wb_clk_i soc.ram_data_out\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_29_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10933_ _05455_ _01371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_204_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10864_ soc.ram_encoder_0.data_out\[6\] _05419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_231_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_220_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10795_ _02223_ soc.spi_video_ram_1.write_fifo.fifo_mem\[7\]\[3\] _05378_ _05382_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XPHY_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_158_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_200_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_185_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_129_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_184_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_199_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_185_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_201_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11416_ _00482_ clknet_leaf_295_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[2\]\[26\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_153_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11347_ _00413_ clknet_leaf_313_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[27\]\[15\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_125_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_165_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11278_ _00344_ clknet_leaf_200_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[1\]\[4\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_106_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10229_ _02237_ soc.spi_video_ram_1.write_fifo.fifo_mem\[5\]\[10\] _05041_ _05042_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_214_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_230_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_227_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5980 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5991 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05770_ soc.ram_data_out\[5\] _01579_ _01573_ net42 _01618_ _01673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_66_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_207_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_223_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07440_ _03021_ soc.spi_video_ram_1.write_fifo.fifo_mem\[19\]\[27\] _02614_ _03089_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_62_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07371_ _02784_ soc.spi_video_ram_1.write_fifo.fifo_mem\[18\]\[11\] _03020_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_50_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_206_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_149_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_241_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09110_ _04285_ _00717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06322_ _02176_ _00039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_176_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09041_ soc.spi_video_ram_1.write_fifo.read_pointer\[0\] soc.spi_video_ram_1.fifo_read_request
+ _04244_ _04246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_06253_ soc.spi_video_ram_1.fifo_in_data\[5\] _02130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_148_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06184_ _01516_ _01546_ _01471_ _02071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_117_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_239_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09943_ soc.ram_encoder_0.input_bits_left\[4\] _04841_ _04845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_217_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_131_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_154_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_225_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xclkbuf_leaf_161_wb_clk_i clknet_5_27_0_wb_clk_i clknet_leaf_161_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_09874_ _04605_ _04761_ _04762_ _04791_ _04792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_219_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4008 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4019 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08825_ _04129_ _00588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_100_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_180_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05968_ soc.video_generator_1.v_count\[2\] _01861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_08756_ soc.spi_video_ram_1.write_fifo.fifo_mem\[24\]\[14\] _04052_ _04087_ _04092_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_72_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_96_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07707_ soc.spi_video_ram_1.write_fifo.fifo_mem\[0\]\[24\] soc.spi_video_ram_1.write_fifo.fifo_mem\[1\]\[24\]
+ soc.spi_video_ram_1.write_fifo.fifo_mem\[2\]\[24\] soc.spi_video_ram_1.write_fifo.fifo_mem\[3\]\[24\]
+ _02679_ _02894_ _03353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_2628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_148_1423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05899_ _01793_ _01794_ _01795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_08687_ soc.spi_video_ram_1.fifo_in_data\[14\] _04052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_54_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1905 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1927 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_199_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07638_ soc.spi_video_ram_1.write_fifo.fifo_mem\[18\]\[14\] soc.spi_video_ram_1.write_fifo.fifo_mem\[19\]\[14\]
+ _02612_ _03284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_1938 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_246_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_213_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1949 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_202_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07569_ _02784_ soc.spi_video_ram_1.write_fifo.fifo_mem\[14\]\[13\] _03215_ _02647_
+ _03216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_70_1506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09308_ _04404_ _00796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_107_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10580_ _01613_ _05261_ _05263_ _01210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_142_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09239_ _04367_ _00764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_10_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12250_ _01278_ clknet_leaf_135_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[31\]\[3\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_68_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11201_ _00267_ clknet_leaf_46_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[11\]\[11\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_107_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_181_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12181_ _01209_ net87 net77 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_102_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_237_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_194_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_1405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_249_wb_clk_i clknet_5_17_0_wb_clk_i clknet_leaf_249_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_68_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11132_ _00198_ clknet_leaf_310_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[14\]\[12\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_123_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_66_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11063_ _00129_ clknet_leaf_224_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[13\]\[1\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_95_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10014_ _04892_ _01015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_131_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_231_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_133_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_209_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_49_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_114_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_236_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3830 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_149_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3841 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3852 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3863 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11965_ _01024_ clknet_leaf_147_wb_clk_i soc.ram_encoder_0.request_address\[2\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3874 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_205_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3885 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3896 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10916_ soc.spi_video_ram_1.write_fifo.fifo_mem\[8\]\[14\] _04052_ _05442_ _05447_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_229_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11896_ _00955_ clknet_leaf_253_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[3\]\[22\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_189_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_1753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10847_ _05409_ _01331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_53_1726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_207_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_201_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10778_ _03344_ _05358_ _05372_ _01299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_40_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_185_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_236_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_141_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_06940_ _02600_ _02601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_45_1243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06871_ _02438_ _02452_ _02540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05822_ _01716_ _01721_ _01722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08610_ _04009_ _00493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09590_ soc.rom_encoder_0.input_buffer\[0\] _04586_ _04553_ _04595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_110_1500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_83_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05753_ soc.ram_data_out\[4\] _01579_ _01573_ net41 _01563_ _01657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_08541_ _02130_ soc.spi_video_ram_1.write_fifo.fifo_mem\[2\]\[5\] _03967_ _03973_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_70_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08472_ _03936_ _00428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05684_ _01591_ _01592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_51_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_184_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07423_ _02922_ soc.spi_video_ram_1.write_fifo.fifo_mem\[9\]\[27\] _03024_ _03072_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_51_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07354_ soc.spi_video_ram_1.write_fifo.fifo_mem\[24\]\[28\] soc.spi_video_ram_1.write_fifo.fifo_mem\[25\]\[28\]
+ soc.spi_video_ram_1.write_fifo.fifo_mem\[26\]\[28\] soc.spi_video_ram_1.write_fifo.fifo_mem\[27\]\[28\]
+ _02644_ _02646_ _03004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_56_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06305_ soc.spi_video_ram_1.fifo_in_address\[6\] _02165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_34_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07285_ _02926_ soc.spi_video_ram_1.write_fifo.fifo_mem\[15\]\[10\] _02838_ _02935_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xcaravel_hack_soc_109 io_oeb[35] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_09024_ _04063_ _04225_ _04236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_164_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06236_ _02114_ _02117_ _02118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_152_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06167_ soc.spi_video_ram_1.read_value\[2\] soc.spi_video_ram_1.read_value\[3\] _01902_
+ _02060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_144_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06098_ _01989_ _01990_ _01991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_137_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09926_ _02481_ _02482_ _04830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_132_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09857_ _04596_ _04761_ _04762_ _04778_ _04779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_213_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3104 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_218_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08808_ _04120_ _00580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_86_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3115 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09788_ _02268_ soc.spi_video_ram_1.write_fifo.fifo_mem\[3\]\[25\] _04696_ _04724_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_73_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3126 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3137 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3148 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3159 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08739_ soc.spi_video_ram_1.write_fifo.fifo_mem\[24\]\[6\] _02403_ _04076_ _04083_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_2436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1702 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_242_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1713 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11750_ _00811_ clknet_leaf_287_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[4\]\[23\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1724 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1735 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1746 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_187_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10701_ _05331_ _01263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_197_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1768 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_241_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11681_ _00742_ clknet_leaf_129_wb_clk_i soc.video_generator_1.v_count\[9\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_2
XTAP_1779 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_230_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_198_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10632_ _05294_ _01231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_167_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10563_ soc.boot_loading_offset\[3\] _05250_ _05252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_6_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_202_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12302_ _01330_ clknet_leaf_295_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[7\]\[26\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_5_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10494_ soc.cpu.PC.REG.data\[11\] _05206_ _05209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_155_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12233_ _01261_ clknet_leaf_312_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[29\]\[15\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_170_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_237_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12164_ _01192_ clknet_leaf_151_wb_clk_i soc.ram_encoder_0.address\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_69_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11115_ _00181_ clknet_leaf_304_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[12\]\[24\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_150_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_12095_ _01123_ net86 soc.cpu.ALU.x\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_122_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11046_ _00112_ clknet_leaf_320_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[0\]\[13\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_5040 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5051 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5062 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_7_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_5073 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5084 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_237_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5095 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_49_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_4361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3693 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11948_ _01007_ clknet_leaf_148_wb_clk_i soc.ram_encoder_0.request_data_out\[1\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_244_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2970 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_232_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2981 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2992 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_127_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11879_ _00938_ clknet_leaf_214_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[3\]\[5\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_127_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_242_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_220_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_186_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_179_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07070_ _02704_ soc.spi_video_ram_1.write_fifo.fifo_mem\[28\]\[2\] _02728_ _02729_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_179_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_161_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06021_ _01910_ _01913_ _01914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_145_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07972_ soc.spi_video_ram_1.write_fifo.fifo_mem\[20\]\[19\] soc.spi_video_ram_1.write_fifo.fifo_mem\[21\]\[19\]
+ soc.spi_video_ram_1.write_fifo.fifo_mem\[22\]\[19\] soc.spi_video_ram_1.write_fifo.fifo_mem\[23\]\[19\]
+ _02681_ _02758_ _03613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_64_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09711_ net58 _04676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_136_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06923_ soc.spi_video_ram_1.write_fifo.fifo_mem\[8\]\[0\] soc.spi_video_ram_1.write_fifo.fifo_mem\[9\]\[0\]
+ soc.spi_video_ram_1.write_fifo.fifo_mem\[10\]\[0\] soc.spi_video_ram_1.write_fifo.fifo_mem\[11\]\[0\]
+ _02575_ _02578_ _02584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_228_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09642_ _04629_ _00906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06854_ _02435_ _02524_ _02525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_151_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05805_ soc.ram_data_out\[7\] _01579_ _01573_ net44 _01618_ _01706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_06785_ _02463_ _02458_ _02464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_09573_ _04579_ _04582_ _00884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_24_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_224_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05736_ soc.cpu.AReg.data\[1\] _01566_ _01641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08524_ _02175_ soc.spi_video_ram_1.write_fifo.fifo_mem\[28\]\[27\] _03933_ _03963_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_58_1445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05667_ _01564_ _01567_ _01572_ _01575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_08455_ _03925_ _00422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_223_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_212_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07406_ soc.spi_video_ram_1.write_fifo.fifo_mem\[0\]\[11\] soc.spi_video_ram_1.write_fifo.fifo_mem\[1\]\[11\]
+ soc.spi_video_ram_1.write_fifo.fifo_mem\[2\]\[11\] soc.spi_video_ram_1.write_fifo.fifo_mem\[3\]\[11\]
+ _03054_ _02690_ _03055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_08386_ soc.spi_video_ram_1.write_fifo.fifo_mem\[26\]\[21\] _02260_ _03865_ _03889_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_196_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05598_ soc.spi_video_ram_1.output_buffer\[17\] _01507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_52_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07337_ _02651_ soc.spi_video_ram_1.write_fifo.fifo_mem\[6\]\[28\] _02690_ _02987_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_143_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07268_ _01387_ _01386_ soc.spi_video_ram_1.state_sram_clk_counter\[0\] _01390_ _02918_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_178_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09007_ _03189_ _04224_ _04227_ _00672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06219_ _02091_ _02103_ _02104_ _02105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_30_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07199_ soc.spi_video_ram_1.write_fifo.fifo_mem\[16\]\[7\] soc.spi_video_ram_1.write_fifo.fifo_mem\[17\]\[7\]
+ soc.spi_video_ram_1.write_fifo.fifo_mem\[18\]\[7\] soc.spi_video_ram_1.write_fifo.fifo_mem\[19\]\[7\]
+ _02769_ _02770_ _02852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_145_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_116_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_82_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_43_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09909_ soc.rom_encoder_0.toggled_sram_sck _02437_ _04818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_232_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_219_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_210_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_150_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11802_ _00862_ clknet_leaf_291_wb_clk_i soc.spi_video_ram_1.fifo_in_address\[5\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_214_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11733_ _00794_ clknet_leaf_245_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[4\]\[6\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_70_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_199_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_70_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_208_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_30_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_243_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_202_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11664_ _00725_ clknet_leaf_66_wb_clk_i soc.spi_video_ram_1.state_counter\[3\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_186_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_161_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10615_ _05285_ _01223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xclkbuf_leaf_264_wb_clk_i clknet_5_6_0_wb_clk_i clknet_leaf_264_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_11595_ _00661_ clknet_leaf_136_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[21\]\[2\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_122_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_128_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10546_ soc.ram_encoder_0.address\[14\] soc.cpu.AReg.data\[14\] _05227_ _05243_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_227_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_10_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_196_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10477_ _04656_ _05193_ _05196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_182_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_68_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12216_ _01244_ clknet_leaf_264_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[19\]\[27\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_83_1516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_155_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12147_ _01175_ net88 soc.cpu.PC.REG.data\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_151_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_123_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12078_ soc.cpu.PC.in\[1\] net85 soc.cpu.AReg.data\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_65_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11029_ _00095_ clknet_leaf_236_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[16\]\[25\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_110_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_37_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_4180 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_206_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06570_ soc.spi_video_ram_1.write_fifo.fifo_mem\[13\]\[9\] _02235_ _02317_ _02327_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_59_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_233_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05521_ _01420_ soc.spi_video_ram_1.state_sram_clk_counter\[1\] _01421_ _01433_ _01434_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_205_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08240_ _02558_ _03800_ _03801_ _00331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_33_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_221_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_15 net44 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08171_ _03751_ _00312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_192_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_222_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07122_ _02744_ soc.spi_video_ram_1.write_fifo.fifo_mem\[6\]\[4\] _02778_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_174_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07053_ _02644_ _02712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_174_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06004_ _01860_ _01863_ _01897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_138_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_153_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5809 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_233_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_25_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_68_wb_clk_i clknet_5_11_0_wb_clk_i clknet_leaf_68_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_07955_ soc.spi_video_ram_1.output_buffer\[5\] _02676_ _03597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_68_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_229_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_214_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06906_ _00004_ _02567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_233_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07886_ _02971_ soc.spi_video_ram_1.write_fifo.fifo_mem\[6\]\[21\] _03528_ _02827_
+ _03529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_09625_ _04620_ _00898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06837_ soc.ram_encoder_0.output_bits_left\[2\] _02494_ _02510_ _02511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_56_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09556_ soc.rom_encoder_0.input_bits_left\[3\] _04568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_43_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_102_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06768_ _02435_ _02433_ _02447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_58_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_70_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08507_ _03954_ _00445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05719_ _01618_ _01619_ _01620_ _01624_ soc.cpu.ALU.zy _01625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_54_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06699_ soc.spi_video_ram_1.write_fifo.fifo_mem\[14\]\[5\] _02401_ _02391_ _02402_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_09487_ _01463_ _04525_ _04528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_246_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08438_ soc.spi_video_ram_1.write_fifo.fifo_mem\[27\]\[16\] _02335_ _03910_ _03917_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_51_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_197_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_1442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_240_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_225_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_211_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_168_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_162_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08369_ _03880_ _00381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_10400_ _02250_ soc.spi_video_ram_1.write_fifo.fifo_mem\[6\]\[16\] _05135_ _05142_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_11380_ _00446_ clknet_leaf_71_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[28\]\[19\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_178_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10331_ soc.cpu.ALU.x\[0\] _05104_ _05105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_109_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_197_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10262_ _03256_ _05044_ _05059_ _01096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_238_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12001_ _01060_ clknet_leaf_163_wb_clk_i soc.ram_encoder_0.initializing_step\[1\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_121_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10193_ soc.hack_clock_0.counter\[2\] _05018_ _05021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_78_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2030 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2041 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2052 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_234_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2063 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_215_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2074 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2085 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2096 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11716_ _00777_ clknet_leaf_25_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[9\]\[18\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_203_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_226_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_174_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_187_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11647_ _00708_ clknet_leaf_308_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[20\]\[15\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_89_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput13 io_in[26] net13 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_122_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_204_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xinput24 la_data_in[15] net24 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput35 la_data_in[25] net35 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_183_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11578_ _00644_ clknet_leaf_8_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[22\]\[14\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_89_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10529_ _05234_ _01188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_109_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_157_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_217_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_217_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_26_1753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_215_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07740_ _02764_ soc.spi_video_ram_1.write_fifo.fifo_mem\[22\]\[15\] _03385_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_133_1171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_238_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07671_ _02581_ _03314_ _03316_ _03317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09410_ soc.rom_encoder_0.request_address\[6\] _02520_ soc.rom_encoder_0.output_buffer\[3\]
+ _04467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_65_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06622_ _02358_ _00157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_80_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_197_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09341_ _04421_ _00812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06553_ _02318_ _00128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_179_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_186_wb_clk_i clknet_5_28_0_wb_clk_i clknet_leaf_186_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_244_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05504_ soc.spi_video_ram_1.current_state\[4\] _01419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
X_09272_ _03537_ _04375_ _04384_ _00780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06484_ _02278_ _02279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
Xclkbuf_leaf_115_wb_clk_i clknet_5_26_0_wb_clk_i clknet_leaf_115_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_08223_ _02503_ _02483_ _03788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_14_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_193_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_140_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08154_ _03742_ _00304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_162_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07105_ _02685_ _02761_ _02720_ _02762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08085_ soc.spi_video_ram_1.write_fifo.fifo_mem\[11\]\[20\] _02343_ _03679_ _03702_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_146_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_1279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07036_ _02694_ _02695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_162_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_192_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4905 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08987_ soc.spi_video_ram_1.write_fifo.fifo_mem\[21\]\[5\] _02401_ _04210_ _04216_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_4916 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4927 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4938 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07938_ _03577_ _03578_ _03579_ _03580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_102_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4949 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_56_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_228_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_186_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07869_ _02764_ soc.spi_video_ram_1.write_fifo.fifo_mem\[14\]\[22\] _03512_ _02958_
+ _03513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_83_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09608_ soc.rom_encoder_0.input_buffer\[10\] _04607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_244_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_189_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10880_ soc.ram_encoder_0.data_out\[14\] _05427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_216_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09539_ _02116_ _04555_ _04254_ _04559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_19_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_223_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_73_1559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_240_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_19_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_199_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_19_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11501_ _00567_ clknet_leaf_298_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[24\]\[24\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_8_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_156_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_169_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_123_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11432_ _00498_ clknet_leaf_311_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[30\]\[13\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_7_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11363_ _00429_ clknet_leaf_258_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[28\]\[2\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10314_ soc.rom_loader.current_address\[11\] _05092_ _05093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_125_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11294_ _00360_ clknet_leaf_44_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[1\]\[20\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_3_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10245_ _02252_ soc.spi_video_ram_1.write_fifo.fifo_mem\[5\]\[17\] _05041_ _05051_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_26_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10176_ _05007_ _05005_ _05008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_234_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_47_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_245_1442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_143_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_230_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_175_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_191_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_239_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_1446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08910_ soc.spi_video_ram_1.write_fifo.fifo_mem\[25\]\[28\] _02353_ _04143_ _04174_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_63_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09890_ _02456_ _02448_ _04614_ _02443_ _04804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XTAP_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_170_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_213_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08841_ _03335_ _04124_ _04137_ _00596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_69_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08772_ soc.spi_video_ram_1.write_fifo.fifo_mem\[24\]\[22\] _04063_ _04075_ _04100_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_85_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05984_ soc.boot_loading_offset\[2\] _01859_ _01864_ _01877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_239_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07723_ _02644_ _03368_ _03369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_113_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_187_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_65_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_226_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07654_ soc.spi_video_ram_1.write_fifo.fifo_mem\[29\]\[14\] _03300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_168_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_240_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06605_ _02347_ _00151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_53_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_179_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07585_ soc.spi_video_ram_1.write_fifo.fifo_mem\[18\]\[25\] soc.spi_video_ram_1.write_fifo.fifo_mem\[19\]\[25\]
+ _02591_ _03232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_55_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09324_ _02250_ soc.spi_video_ram_1.write_fifo.fifo_mem\[4\]\[16\] _04406_ _04413_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06536_ _02171_ soc.spi_video_ram_1.write_fifo.fifo_mem\[0\]\[25\] _02278_ _02306_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_222_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09255_ _04050_ _04375_ _04376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_55_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_181_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06467_ soc.spi_video_ram_1.write_fifo.fifo_mem\[16\]\[24\] _02266_ _02216_ _02267_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_08206_ soc.rom_encoder_0.initializing_step\[4\] soc.rom_encoder_0.initializing_step\[3\]
+ _02452_ _03775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_09186_ _01853_ _04336_ _04337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06398_ _02220_ _00071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_88_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_1524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08137_ _02122_ soc.spi_video_ram_1.write_fifo.fifo_mem\[10\]\[1\] _03732_ _03734_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_179_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_218_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_190_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_83_wb_clk_i clknet_5_10_0_wb_clk_i clknet_leaf_83_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_200_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08068_ _03693_ _00267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_150_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6104 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_12_wb_clk_i clknet_5_2_0_wb_clk_i clknet_leaf_12_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_07019_ _02643_ _02678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_6115 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6126 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6137 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6148 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10030_ soc.ram_encoder_0.request_address\[1\] soc.ram_encoder_0.address\[1\] _04900_
+ _04901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_5414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6159 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_7_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_5425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_235_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_5447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4702 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4713 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4724 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4735 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4746 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4757 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4768 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_229_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4779 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11981_ _01040_ clknet_leaf_156_wb_clk_i soc.ram_data_out\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_17_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_229_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_232_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10932_ soc.spi_video_ram_1.write_fifo.fifo_mem\[8\]\[22\] _04063_ _05430_ _05455_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_84_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_245_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10863_ _01680_ _05222_ _05412_ _05418_ _01338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_147_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_38_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_34_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10794_ _05381_ _01306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_160_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_185_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_212_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_157_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_16_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_240_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_200_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11415_ _00481_ clknet_leaf_229_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[2\]\[25\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_158_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11346_ _00412_ clknet_leaf_318_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[27\]\[14\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_193_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11277_ _00343_ clknet_leaf_259_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[1\]\[3\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_171_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_239_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10228_ _05029_ _05041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_67_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10159_ _02482_ _04993_ _04553_ _04996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_121_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5970 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_181_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5981 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5992 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_23_1756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_208_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_169_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_165_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_222_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07370_ _02918_ _03019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_210_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_204_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_176_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06321_ _02175_ soc.spi_video_ram_1.write_fifo.fifo_mem\[18\]\[27\] _02119_ _02176_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_143_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09040_ soc.spi_video_ram_1.fifo_read_request _04244_ soc.spi_video_ram_1.write_fifo.read_pointer\[0\]
+ _04245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06252_ _02129_ _00016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_198_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06183_ _01857_ _02070_ net74 vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_30_1749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_190_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_219_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09942_ soc.ram_encoder_0.input_bits_left\[4\] _04841_ _04844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_48_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09873_ soc.rom_encoder_0.request_data_out\[13\] _04742_ _04791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_135_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4009 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08824_ _02153_ soc.spi_video_ram_1.write_fifo.fifo_mem\[23\]\[16\] _04117_ _04129_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_97_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_246_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08755_ _04091_ _00556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_85_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05967_ soc.video_generator_1.v_count\[9\] _01860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_3
XFILLER_22_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_230_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07706_ _03334_ _03342_ _03351_ _00004_ _03352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_2618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_214_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_241_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_227_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08686_ _03214_ _04046_ _04051_ _00527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xclkbuf_leaf_130_wb_clk_i clknet_5_13_0_wb_clk_i clknet_leaf_130_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_05898_ _01756_ _01789_ _01794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_1906 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_241_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_198_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1917 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07637_ soc.video_generator_1.v_count\[3\] _01897_ _03283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_1928 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1939 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_224_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07568_ _02712_ _03214_ _03215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_167_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09307_ _02233_ soc.spi_video_ram_1.write_fifo.fifo_mem\[4\]\[8\] _04395_ _04404_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_55_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06519_ _02297_ _00115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_139_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_194_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07499_ soc.spi_video_ram_1.write_fifo.fifo_mem\[16\]\[26\] soc.spi_video_ram_1.write_fifo.fifo_mem\[17\]\[26\]
+ soc.spi_video_ram_1.write_fifo.fifo_mem\[18\]\[26\] soc.spi_video_ram_1.write_fifo.fifo_mem\[19\]\[26\]
+ _02907_ _02908_ _03147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_16_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09238_ _02227_ soc.spi_video_ram_1.write_fifo.fifo_mem\[9\]\[5\] _04365_ _04367_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_33_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_182_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09169_ _04317_ _04324_ _04325_ _00736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_182_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_237_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_11200_ _00266_ clknet_leaf_15_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[11\]\[10\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_159_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_12180_ _01208_ clknet_leaf_127_wb_clk_i soc.hack_wait_clocks\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_135_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_1447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_190_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_190_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_1428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11131_ _00197_ clknet_leaf_46_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[14\]\[11\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_122_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11062_ _00128_ clknet_leaf_177_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[13\]\[0\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_5211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_88_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_289_wb_clk_i clknet_5_5_0_wb_clk_i clknet_leaf_289_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_237_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10013_ soc.ram_encoder_0.request_data_out\[9\] soc.ram_encoder_0.data_out\[9\] _04889_
+ _04892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_5244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_218_wb_clk_i clknet_5_21_0_wb_clk_i clknet_leaf_218_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_5266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3820 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_4576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3831 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3842 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3853 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_151_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11964_ _01023_ clknet_leaf_149_wb_clk_i soc.ram_encoder_0.request_address\[1\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3864 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_233_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_204_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3875 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3886 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3897 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10915_ _05446_ _01362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_72_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11895_ _00954_ clknet_leaf_230_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[3\]\[21\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_60_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_220_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10846_ _02272_ soc.spi_video_ram_1.write_fifo.fifo_mem\[7\]\[27\] _05389_ _05409_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_34_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10777_ _04067_ _05359_ _05372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_12_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_199_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_201_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_1484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_12_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_172_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11329_ _00395_ clknet_leaf_292_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[26\]\[26\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_119_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_214_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06870_ _02528_ _01592_ _02539_ _01555_ _00224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_68_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_171_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_227_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05821_ _01705_ _01720_ _01721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_10_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_114_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08540_ _03972_ _00460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_78_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05752_ _01557_ _01655_ _01656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_209_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_223_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_93_1529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08471_ _02122_ soc.spi_video_ram_1.write_fifo.fifo_mem\[28\]\[1\] _03934_ _03936_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_05683_ soc.cpu.instruction\[15\] _01590_ _01591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_243_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07422_ _02971_ soc.spi_video_ram_1.write_fifo.fifo_mem\[8\]\[27\] _03071_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_196_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_165_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_225_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_211_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_206_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_149_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07353_ _02601_ _03002_ _03003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_176_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06304_ _02164_ _00033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_108_1496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07284_ _02924_ soc.spi_video_ram_1.write_fifo.fifo_mem\[14\]\[10\] _02934_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_108_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09023_ _03557_ _04224_ _04235_ _00680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06235_ _02115_ _01403_ _02116_ _02117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_102_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_191_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06166_ _01839_ _01846_ _02059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_132_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_191_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06097_ soc.video_generator_1.h_count\[1\] soc.display_clks_before_active\[0\] _01990_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_132_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09925_ _04787_ soc.ram_encoder_0.toggled_sram_sck _00989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_120_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_219_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09856_ soc.rom_encoder_0.request_data_out\[9\] _04742_ _04778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_311_wb_clk_i clknet_5_1_0_wb_clk_i clknet_leaf_311_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_100_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08807_ _02136_ soc.spi_video_ram_1.write_fifo.fifo_mem\[23\]\[8\] _04117_ _04120_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_98_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3105 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09787_ _04723_ _00957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3116 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_189_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06999_ _02596_ _02658_ _02659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_3127 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3138 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3149 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08738_ _04082_ _00548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_215_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_199_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1714 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1725 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08669_ _04040_ _00521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_42_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1736 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_202_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1747 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10700_ _02252_ soc.spi_video_ram_1.write_fifo.fifo_mem\[29\]\[17\] _05321_ _05331_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_148_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1769 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11680_ _00741_ clknet_leaf_63_wb_clk_i soc.video_generator_1.v_count\[8\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_183_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_243_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_201_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10631_ soc.spi_video_ram_1.write_fifo.fifo_mem\[19\]\[14\] _04052_ _05289_ _05294_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_70_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_204_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_197_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_220_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10562_ soc.boot_loading_offset\[3\] _05250_ _05251_ _01204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_126_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12301_ _01329_ clknet_leaf_289_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[7\]\[25\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_127_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_212_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_196_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_182_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10493_ _05172_ _05207_ _05208_ _01177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_6_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12232_ _01260_ clknet_leaf_316_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[29\]\[14\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_107_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12163_ _01191_ clknet_leaf_148_wb_clk_i soc.ram_encoder_0.address\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_29_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11114_ _00180_ clknet_leaf_236_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[12\]\[23\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_81_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12094_ _01122_ net86 soc.cpu.ALU.x\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_89_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5030 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11045_ _00111_ clknet_leaf_0_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[0\]\[12\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_231_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5041 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5052 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_1488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_209_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5063 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5074 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5085 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5096 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_205_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11947_ _01006_ clknet_leaf_152_wb_clk_i soc.ram_encoder_0.request_data_out\[0\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_73_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_1384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3694 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_229_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2960 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2971 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_221_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_189_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_178_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2982 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2993 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11878_ _00937_ clknet_leaf_199_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[3\]\[4\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_207_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10829_ _05400_ _01322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_32_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_186_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_186_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_125_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06020_ _01844_ _01912_ _01913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_127_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_47_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_236_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07971_ _02768_ _03611_ _03612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_68_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09710_ _04675_ _00928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06922_ _02582_ _02583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_132_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09641_ soc.rom_encoder_0.data_out\[8\] soc.rom_encoder_0.request_data_out\[8\] _04621_
+ _04629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06853_ _02434_ _02454_ _02524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_99_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_3_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05804_ _01561_ _01705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_132_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09572_ soc.rom_encoder_0.input_bits_left\[4\] _04580_ _04582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_110_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06784_ _02462_ _02463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_71_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08523_ _03962_ _00453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05735_ net40 _01640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_36_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_227_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_184_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08454_ soc.spi_video_ram_1.write_fifo.fifo_mem\[27\]\[24\] _02266_ _03898_ _03925_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_51_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05666_ net29 _01573_ _01574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07405_ _02902_ _03054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_11_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_56_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08385_ _03888_ _00389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_123_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05597_ _01486_ _01502_ _01505_ _01506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_177_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07336_ _02941_ soc.spi_video_ram_1.write_fifo.fifo_mem\[7\]\[28\] _02986_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_221_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07267_ _02055_ _02916_ _02917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_136_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09006_ _04050_ _04225_ _04227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_139_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06218_ _01492_ _01484_ _02104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07198_ soc.spi_video_ram_1.write_fifo.fifo_mem\[20\]\[7\] soc.spi_video_ram_1.write_fifo.fifo_mem\[21\]\[7\]
+ soc.spi_video_ram_1.write_fifo.fifo_mem\[22\]\[7\] soc.spi_video_ram_1.write_fifo.fifo_mem\[23\]\[7\]
+ _02764_ _02723_ _02851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_121_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_195_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_1406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06149_ _02027_ _02029_ _02030_ _01864_ _02041_ _02042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_105_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_219_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09908_ _02459_ _04731_ soc.rom_encoder_0.initializing_step\[1\] _04817_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_150_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_101_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09839_ _04752_ _04765_ _00967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_246_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_210_1753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_234_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11801_ _00861_ clknet_leaf_55_wb_clk_i soc.spi_video_ram_1.fifo_in_address\[4\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_162_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_3_1_0_wb_clk_i clknet_2_0_0_wb_clk_i clknet_3_1_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_55_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_26_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_203_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11732_ _00793_ clknet_leaf_227_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[4\]\[5\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_226_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_2289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_230_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_11663_ _00724_ clknet_leaf_65_wb_clk_i soc.spi_video_ram_1.state_counter\[2\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_14_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10614_ soc.spi_video_ram_1.write_fifo.fifo_mem\[19\]\[6\] _02403_ _05278_ _05285_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_168_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11594_ _00660_ clknet_leaf_208_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[21\]\[1\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10545_ _01456_ _05228_ _05242_ _01196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_183_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_155_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10476_ _05171_ _05194_ _05195_ _01173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_155_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12215_ _01243_ clknet_leaf_288_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[19\]\[26\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_237_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_233_wb_clk_i clknet_5_5_0_wb_clk_i clknet_leaf_233_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_100_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_174_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12146_ _01174_ net89 soc.cpu.PC.REG.data\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_123_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_238_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12077_ soc.cpu.PC.in\[0\] net84 soc.cpu.AReg.data\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_42_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11028_ _00094_ clknet_leaf_304_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[16\]\[24\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_65_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_237_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4170 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4181 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_244_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05520_ _01432_ soc.spi_video_ram_1.state_sram_clk_counter\[6\] soc.spi_video_ram_1.state_sram_clk_counter\[5\]
+ soc.spi_video_ram_1.state_sram_clk_counter\[4\] _01433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_166_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_146_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2790 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_127_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_220_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_16 net78 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_159_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08170_ _02155_ soc.spi_video_ram_1.write_fifo.fifo_mem\[10\]\[17\] _03743_ _03751_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_105_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_140_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07121_ _02697_ soc.spi_video_ram_1.write_fifo.fifo_mem\[5\]\[4\] _02742_ _02777_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_203_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_146_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07052_ _02684_ _02687_ _02709_ _02710_ _02711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_06003_ _01852_ _01854_ _01857_ _01867_ _01896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_192_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_130_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_141_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07954_ _02677_ _01392_ _02734_ _03596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_228_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06905_ _02556_ _02565_ _02566_ _00232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07885_ _02688_ _03527_ _03528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_99_1535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_151_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09624_ soc.rom_encoder_0.data_out\[0\] soc.rom_encoder_0.request_data_out\[0\] _04618_
+ _04620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_83_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_216_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06836_ _02482_ _02497_ _02510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_09555_ soc.rom_encoder_0.current_state\[2\] _02447_ _04567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_243_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06767_ soc.rom_encoder_0.request_write _02443_ _02445_ _02446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
Xclkbuf_leaf_37_wb_clk_i clknet_5_3_0_wb_clk_i clknet_leaf_37_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_97_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08506_ _02157_ soc.spi_video_ram_1.write_fifo.fifo_mem\[28\]\[18\] _03945_ _03954_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_05718_ _01573_ _01621_ _01622_ _01623_ _01624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_09486_ _04519_ _04525_ _04527_ _00852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_227_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06698_ soc.spi_video_ram_1.fifo_in_data\[5\] _02401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_212_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08437_ _03916_ _00413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_169_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05649_ soc.cpu.ALU.nx _01557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_196_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08368_ soc.spi_video_ram_1.write_fifo.fifo_mem\[26\]\[12\] _02242_ _03877_ _03880_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_240_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07319_ _02620_ _02947_ _02968_ _02969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_20_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08299_ _03829_ _03842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_137_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_194_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10330_ _05102_ _05104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_192_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10261_ soc.spi_video_ram_1.fifo_in_address\[9\] _05045_ _05059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_12000_ _01059_ clknet_leaf_163_wb_clk_i soc.ram_encoder_0.initializing_step\[0\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_106_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_234_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10192_ soc.hack_clock_0.counter\[2\] _05018_ _05020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_156_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_191_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_232_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_219_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_235_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_185_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2020 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2031 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2042 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2053 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2064 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2075 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2086 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_167_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2097 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_199_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11715_ _00776_ clknet_leaf_24_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[9\]\[17\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_202_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11646_ _00707_ clknet_leaf_6_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[20\]\[14\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xinput14 io_in[30] net14 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
Xinput25 la_data_in[16] net25 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_128_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_156_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput36 la_data_in[26] net36 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_11577_ _00643_ clknet_leaf_40_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[22\]\[13\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_141_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10528_ soc.ram_encoder_0.address\[5\] soc.cpu.AReg.data\[5\] _05227_ _05234_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_156_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_196_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10459_ _05171_ _05181_ _05182_ _01169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_124_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12129_ _01157_ clknet_leaf_289_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[6\]\[21\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_112_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07670_ _02695_ soc.spi_video_ram_1.write_fifo.fifo_mem\[13\]\[14\] _03315_ _02741_
+ _03316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_93_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_203_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06621_ _02113_ soc.spi_video_ram_1.write_fifo.fifo_mem\[12\]\[0\] _02357_ _02358_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_225_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_1279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09340_ _02266_ soc.spi_video_ram_1.write_fifo.fifo_mem\[4\]\[24\] _04394_ _04421_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_94_1443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06552_ soc.spi_video_ram_1.write_fifo.fifo_mem\[13\]\[0\] _02310_ _02317_ _02318_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_80_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05503_ _01409_ _01417_ _01418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_09271_ _04061_ _04360_ _04384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_61_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06483_ _02277_ _02278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_221_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_33_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08222_ _02556_ _03786_ _03787_ _00327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_146_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_222_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08153_ _02138_ soc.spi_video_ram_1.write_fifo.fifo_mem\[10\]\[9\] _03732_ _03742_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_147_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_155_wb_clk_i clknet_5_30_0_wb_clk_i clknet_leaf_155_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_101_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_147_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07104_ soc.spi_video_ram_1.write_fifo.fifo_mem\[20\]\[3\] soc.spi_video_ram_1.write_fifo.fifo_mem\[21\]\[3\]
+ soc.spi_video_ram_1.write_fifo.fifo_mem\[22\]\[3\] soc.spi_video_ram_1.write_fifo.fifo_mem\[23\]\[3\]
+ _02717_ _02682_ _02761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_119_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_200_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_174_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08084_ _03701_ _00275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_101_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07035_ _02572_ _02694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_162_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_114_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_5607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_103_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08986_ _04215_ _00663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_103_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_233_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4906 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4917 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_229_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4928 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07937_ _02831_ _03579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_112_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4939 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07868_ _02635_ _03511_ _03512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_217_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06819_ soc.ram_encoder_0.output_bits_left\[3\] _02494_ _02495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09607_ _04605_ _04585_ _04606_ _00894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_3_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07799_ _03054_ _03443_ _03444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_186_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09538_ _01446_ _04552_ _04558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XPHY_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_184_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_12_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09469_ _02443_ _04513_ _04514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XPHY_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_125_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_197_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11500_ _00566_ clknet_leaf_234_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[24\]\[23\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_240_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_200_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_178_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_8_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11431_ _00497_ clknet_leaf_6_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[30\]\[12\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_125_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11362_ _00428_ clknet_leaf_224_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[28\]\[1\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_193_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_197_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10313_ _05071_ _05091_ _05092_ _01113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_98_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11293_ _00359_ clknet_leaf_68_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[1\]\[19\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_238_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_5_22_0_wb_clk_i clknet_4_11_0_wb_clk_i clknet_5_22_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_10244_ _05050_ _01087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_152_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_133_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10175_ soc.ram_encoder_0.initializing_step\[3\] _05007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_117_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_212_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_207_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_234_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_76_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_31_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1171 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_203_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_188_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_176_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_187_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11629_ _00007_ clknet_leaf_69_wb_clk_i soc.spi_video_ram_1.current_state\[2\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_204_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_184_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08840_ _04067_ _04110_ _04137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_44_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08771_ _04099_ _00564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_230_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_215_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05983_ _01858_ _01865_ _01868_ _01875_ _01876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_4
XTAP_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_245_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_238_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07722_ soc.spi_video_ram_1.write_fifo.fifo_mem\[15\]\[24\] _03368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_6_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07653_ _02574_ soc.spi_video_ram_1.write_fifo.fifo_mem\[30\]\[14\] _03298_ _02894_
+ _03299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_26_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06604_ soc.spi_video_ram_1.write_fifo.fifo_mem\[13\]\[23\] _02264_ _02316_ _02347_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_187_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07584_ _02710_ _03207_ _03230_ _03019_ _03231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_41_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_228_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09323_ _04412_ _00803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_179_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06535_ _02305_ _00123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_240_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_181_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09254_ _04359_ _04375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_06466_ soc.spi_video_ram_1.fifo_in_address\[8\] _02266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_22_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_193_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08205_ _03763_ _02449_ _03773_ _03774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_21_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_194_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09185_ _04317_ _04335_ _04336_ _00741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_239_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06397_ soc.spi_video_ram_1.write_fifo.fifo_mem\[16\]\[1\] _02219_ _02217_ _02220_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_147_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08136_ _03733_ _00295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_175_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_162_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_190_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_179_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08067_ soc.spi_video_ram_1.write_fifo.fifo_mem\[11\]\[11\] _02414_ _03691_ _03693_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_135_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07018_ soc.spi_video_ram_1.current_state\[1\] _02677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_6105 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_162_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6116 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_89_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6127 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6138 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6149 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_192_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_88_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_216_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4703 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4714 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xclkbuf_leaf_52_wb_clk_i clknet_5_13_0_wb_clk_i clknet_leaf_52_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_4725 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_170_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08969_ soc.spi_video_ram_1.write_fifo.fifo_mem\[22\]\[26\] _03927_ _04177_ _04206_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_130_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4736 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4747 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4758 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11980_ _01039_ clknet_leaf_157_wb_clk_i soc.ram_data_out\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_4769 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10931_ _05454_ _01370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_79_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_244_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_216_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10862_ soc.ram_encoder_0.data_out\[5\] _05418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_147_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_1752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_207_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_232_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_77_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_242_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_73_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10793_ _02221_ soc.spi_video_ram_1.write_fifo.fifo_mem\[7\]\[2\] _05378_ _05381_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XPHY_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_207_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_33_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_205_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_166_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11414_ _00480_ clknet_leaf_299_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[2\]\[24\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_51_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_165_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11345_ _00411_ clknet_leaf_315_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[27\]\[13\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_181_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11276_ _00342_ clknet_leaf_258_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[1\]\[2\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_136_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10227_ _05040_ _01080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_234_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10158_ soc.ram_encoder_0.request_write _04831_ _04874_ _04994_ _04995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_67_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_239_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5960 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5971 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_5982 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5993 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10089_ soc.ram_data_out\[2\] _04927_ _04941_ _04942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_236_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_235_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_245_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_200_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_222_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06320_ soc.spi_video_ram_1.fifo_in_address\[11\] _02175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_176_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_06251_ _02128_ soc.spi_video_ram_1.write_fifo.fifo_mem\[18\]\[4\] _02120_ _02129_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_191_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06182_ _01853_ _01931_ soc.video_generator_1.v_count\[2\] _02069_ _02070_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_102_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09941_ _04841_ _04842_ _04843_ _00991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_132_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_213_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09872_ _04787_ _04790_ _00975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_1559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08823_ _04128_ _00587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_189_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_85_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_239_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08754_ soc.spi_video_ram_1.write_fifo.fifo_mem\[24\]\[13\] _04050_ _04087_ _04091_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_61_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05966_ soc.video_generator_1.v_count\[9\] _01850_ _01851_ _01859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_113_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07705_ _02706_ _03343_ _03350_ _00003_ _03351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_2608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08685_ _04050_ _04048_ _04051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_66_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_226_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05897_ _01792_ _01776_ _01775_ _01793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_54_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1907 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1918 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07636_ _03282_ _00246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_246_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1929 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_214_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07567_ soc.spi_video_ram_1.write_fifo.fifo_mem\[15\]\[13\] _03214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xclkbuf_leaf_170_wb_clk_i clknet_5_31_0_wb_clk_i clknet_leaf_170_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_110_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_241_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09306_ _04403_ _00795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06518_ _02153_ soc.spi_video_ram_1.write_fifo.fifo_mem\[0\]\[16\] _02290_ _02297_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_142_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07498_ _02620_ _03126_ _03145_ _02918_ _03146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_107_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_224_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09237_ _04366_ _00763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06449_ soc.spi_video_ram_1.write_fifo.fifo_mem\[16\]\[18\] _02254_ _02238_ _02255_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_210_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_194_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09168_ soc.video_generator_1.v_count\[3\] _04323_ _04325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_108_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_147_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08119_ _03713_ _03721_ _00290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_120_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_198_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09099_ _02256_ soc.spi_video_ram_1.write_fifo.fifo_mem\[20\]\[19\] _04270_ _04280_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_123_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_163_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11130_ _00196_ clknet_leaf_16_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[14\]\[10\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_123_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_135_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11061_ _00127_ clknet_leaf_296_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[0\]\[28\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_118_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_235_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_77_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_5223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10012_ _04891_ _01014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_5234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_133_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_5245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_5256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_192_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_4511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_4522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_130_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3810 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_218_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3821 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3832 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_229_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3843 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11963_ _01022_ clknet_leaf_148_wb_clk_i soc.ram_encoder_0.request_address\[0\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3854 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3865 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xclkbuf_leaf_258_wb_clk_i clknet_5_18_0_wb_clk_i clknet_leaf_258_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_3876 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3887 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_217_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10914_ soc.spi_video_ram_1.write_fifo.fifo_mem\[8\]\[13\] _04050_ _05442_ _05446_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_3898 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11894_ _00953_ clknet_leaf_45_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[3\]\[20\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_233_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10845_ _03175_ _05392_ _05408_ _01330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_38_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_204_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_198_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_242_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10776_ _03440_ _05358_ _05371_ _01298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_9_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_203_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_240_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_200_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_177_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_1548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_126_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11328_ _00394_ clknet_leaf_231_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[26\]\[25\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_140_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11259_ _00325_ clknet_leaf_149_wb_clk_i soc.ram_encoder_0.output_buffer\[5\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_6480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_80_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_171_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_39_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05820_ _01717_ _01719_ _01720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_94_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5790 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_1502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_243_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05751_ _01558_ soc.cpu.ALU.x\[4\] _01655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_208_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08470_ _03935_ _00427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05682_ soc.cpu.instruction\[5\] _01590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_35_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_208_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_211_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07421_ _03021_ soc.spi_video_ram_1.write_fifo.fifo_mem\[11\]\[27\] _02652_ _03070_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_56_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_210_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_223_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07352_ _02998_ _02999_ _03001_ _02598_ _02900_ _03002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_143_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_188_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06303_ _02163_ soc.spi_video_ram_1.write_fifo.fifo_mem\[18\]\[21\] _02119_ _02164_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_91_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_225_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07283_ _02922_ soc.spi_video_ram_1.write_fifo.fifo_mem\[12\]\[10\] _02932_ _02933_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_149_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09022_ _04061_ _04225_ _04235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06234_ soc.spi_video_ram_1.write_fifo.write_pointer\[2\] _02116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_176_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_129_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_4_3_0_wb_clk_i clknet_3_1_0_wb_clk_i clknet_4_3_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_117_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06165_ _02054_ _02057_ _02058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_219_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_1749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06096_ _01902_ _01903_ _01989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_132_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_176_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09924_ soc.rom_encoder_0.initializing_step\[4\] _04828_ _04829_ _03714_ _00988_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_28_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09855_ _04752_ _04777_ _00971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08806_ _04119_ _00579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_22_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3106 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09786_ _02266_ soc.spi_video_ram_1.write_fifo.fifo_mem\[3\]\[24\] _04696_ _04723_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06998_ soc.spi_video_ram_1.write_fifo.fifo_mem\[28\]\[1\] soc.spi_video_ram_1.write_fifo.fifo_mem\[29\]\[1\]
+ soc.spi_video_ram_1.write_fifo.fifo_mem\[30\]\[1\] soc.spi_video_ram_1.write_fifo.fifo_mem\[31\]\[1\]
+ _02635_ _02636_ _02658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_22_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3117 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_67_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3128 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_230_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3139 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_233_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05949_ _01837_ _01839_ _01842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XTAP_2405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08737_ soc.spi_video_ram_1.write_fifo.fifo_mem\[24\]\[5\] _02401_ _04076_ _04082_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_2416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_227_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_22_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_198_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1704 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08668_ soc.spi_video_ram_1.write_fifo.fifo_mem\[15\]\[7\] _02405_ _04032_ _04040_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_1715 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_183_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_148_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1726 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1737 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_215_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_183_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07619_ soc.spi_video_ram_1.write_fifo.fifo_mem\[9\]\[25\] _03266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_1748 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1759 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08599_ _02126_ soc.spi_video_ram_1.write_fifo.fifo_mem\[30\]\[3\] _04000_ _04004_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_39_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_1411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10630_ _05293_ _01230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_161_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10561_ soc.boot_loading_offset\[3\] _05250_ _04248_ _05251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_10_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12300_ _01328_ clknet_leaf_300_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[7\]\[24\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_6_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_241_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10492_ soc.cpu.PC.in\[11\] _05188_ _05201_ _05208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_136_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12231_ _01259_ clknet_leaf_311_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[29\]\[13\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_205_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12162_ _01190_ clknet_leaf_146_wb_clk_i soc.ram_encoder_0.address\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_122_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11113_ _00179_ clknet_leaf_267_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[12\]\[22\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12093_ _01121_ net86 soc.cpu.ALU.x\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_110_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5020 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11044_ _00110_ clknet_leaf_36_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[0\]\[11\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_104_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5031 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5042 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5053 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_133_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5064 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5075 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5086 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_225_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5097 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11946_ _01005_ clknet_leaf_154_wb_clk_i soc.ram_encoder_0.request_write vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_2_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_209_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2950 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3695 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2961 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2972 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_72_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2983 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11877_ _00936_ clknet_leaf_259_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[3\]\[3\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2994 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_205_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10828_ _02254_ soc.spi_video_ram_1.write_fifo.fifo_mem\[7\]\[18\] _05389_ _05400_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_186_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_199_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10759_ _04054_ _05359_ _05363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_158_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_145_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_220_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_141_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_173_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07970_ soc.spi_video_ram_1.write_fifo.fifo_mem\[16\]\[19\] soc.spi_video_ram_1.write_fifo.fifo_mem\[17\]\[19\]
+ soc.spi_video_ram_1.write_fifo.fifo_mem\[18\]\[19\] soc.spi_video_ram_1.write_fifo.fifo_mem\[19\]\[19\]
+ _02769_ _02770_ _03611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_142_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_214_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06921_ _02581_ _02582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_171_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_06852_ _02513_ _02522_ _02523_ _00222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09640_ _04628_ _00905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_132_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_109_wb_clk_i clknet_5_15_0_wb_clk_i clknet_leaf_109_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_23_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05803_ _01702_ _01703_ _01704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_09571_ _04579_ _04580_ _04581_ _00883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_132_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_215_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06783_ soc.rom_encoder_0.output_bits_left\[4\] _02440_ _02462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_209_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08522_ _02173_ soc.spi_video_ram_1.write_fifo.fifo_mem\[28\]\[26\] _03933_ _03962_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_05734_ _01598_ _01638_ _01639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_58_1414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_70_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_227_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_63_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08453_ _03924_ _00421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05665_ soc.cpu.AReg.data\[0\] _01567_ _01572_ _01573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_51_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_196_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_180_1319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_211_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07404_ _02640_ _03052_ _03053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_36_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08384_ soc.spi_video_ram_1.write_fifo.fifo_mem\[26\]\[20\] _02343_ _03865_ _03888_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_05596_ _01473_ _01504_ _01505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_195_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07335_ soc.spi_video_ram_1.write_fifo.fifo_mem\[0\]\[28\] soc.spi_video_ram_1.write_fifo.fifo_mem\[1\]\[28\]
+ soc.spi_video_ram_1.write_fifo.fifo_mem\[2\]\[28\] soc.spi_video_ram_1.write_fifo.fifo_mem\[3\]\[28\]
+ _02931_ _02690_ _02985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_137_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07266_ _02056_ _02916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09005_ _03112_ _04224_ _04226_ _00671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06217_ _01486_ _01483_ _02103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_118_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_191_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07197_ soc.spi_video_ram_1.write_fifo.fifo_mem\[24\]\[7\] soc.spi_video_ram_1.write_fifo.fifo_mem\[25\]\[7\]
+ soc.spi_video_ram_1.write_fifo.fifo_mem\[26\]\[7\] soc.spi_video_ram_1.write_fifo.fifo_mem\[27\]\[7\]
+ _02769_ _02770_ _02850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_133_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06148_ _01947_ _02033_ _02040_ _01932_ _02041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_133_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_191_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06079_ _01925_ _01971_ _01972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_120_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_236_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09907_ _04816_ _00984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_43_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_76_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09838_ soc.cpu.instruction\[4\] _04740_ _04764_ _04765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_98_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_207_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09769_ _04714_ _00948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11800_ _00860_ clknet_leaf_67_wb_clk_i soc.spi_video_ram_1.fifo_in_address\[3\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_199_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_2257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11731_ _00792_ clknet_leaf_262_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[4\]\[4\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_155_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_187_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_70_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11662_ _00723_ clknet_leaf_64_wb_clk_i soc.spi_video_ram_1.state_counter\[1\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_70_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_204_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10613_ _05284_ _01222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_11593_ _00659_ clknet_leaf_205_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[21\]\[0\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_126_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10544_ soc.ram_encoder_0.address\[13\] _05228_ _05242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_127_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_183_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_196_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_182_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_41_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10475_ soc.cpu.PC.in\[7\] _05188_ _05173_ _05195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_87_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_170_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12214_ _01242_ clknet_leaf_234_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[19\]\[25\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_100_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_83_1518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_233_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_12145_ _01173_ net88 soc.cpu.PC.REG.data\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_2_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_7_wb_clk_i clknet_5_2_0_wb_clk_i clknet_leaf_7_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_69_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_215_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12076_ _01119_ clknet_leaf_129_wb_clk_i net83 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_133_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_273_wb_clk_i clknet_5_6_0_wb_clk_i clknet_leaf_273_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_2_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11027_ _00093_ clknet_leaf_236_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[16\]\[23\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_65_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_202_wb_clk_i clknet_5_19_0_wb_clk_i clknet_leaf_202_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_238_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4160 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4171 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4182 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_52_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_221_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_178_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11929_ _00988_ clknet_leaf_86_wb_clk_i soc.rom_encoder_0.initializing_step\[4\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XTAP_2780 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_181_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2791 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_162_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_242_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07120_ _02726_ soc.spi_video_ram_1.write_fifo.fifo_mem\[4\]\[4\] _02776_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_70_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_179_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07051_ _02655_ _02710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_173_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06002_ soc.boot_loading_offset\[0\] _01895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_115_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_192_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07953_ _03585_ _03594_ _03595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_64_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06904_ soc.ram_encoder_0.output_buffer\[1\] _02563_ _02566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_56_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07884_ soc.spi_video_ram_1.write_fifo.fifo_mem\[7\]\[21\] _03527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_210_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_244_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09623_ _04426_ _04618_ _04619_ _00897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_56_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06835_ _02494_ _02508_ _02509_ _00219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_186_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09554_ _02434_ _02457_ _04566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_06766_ _02433_ _02444_ _02445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_55_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05717_ soc.cpu.AReg.data\[0\] net39 _01567_ _01572_ _01623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or4_1
XFILLER_58_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08505_ _03953_ _00444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_19_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06697_ _02400_ _00190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09485_ _01470_ _04526_ _04527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_197_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_169_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05648_ soc.cpu.ALU.no _01556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_08436_ soc.spi_video_ram_1.write_fifo.fifo_mem\[27\]\[15\] _02248_ _03910_ _03916_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_51_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_77_wb_clk_i clknet_5_8_0_wb_clk_i clknet_leaf_77_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_71_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08367_ _03879_ _00380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05579_ _01463_ _01487_ _01488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_221_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07318_ _02953_ _02960_ _00004_ _02967_ _02968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_109_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_164_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08298_ _03841_ _00349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_197_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07249_ _00002_ _02900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_121_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10260_ _03357_ _05044_ _05058_ _01095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_30_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_5_12_0_wb_clk_i clknet_4_6_0_wb_clk_i clknet_5_12_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_69_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_219_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10191_ _05017_ _05018_ _05019_ _01065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_105_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_121_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_238_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_246_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_234_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_185_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2010 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2021 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2032 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2043 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2054 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2065 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_203_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_226_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2076 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2087 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2098 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_230_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11714_ _00775_ clknet_leaf_76_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[9\]\[16\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_159_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11645_ _00706_ clknet_leaf_39_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[20\]\[13\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_35_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xinput15 io_in[31] net15 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_11576_ _00642_ clknet_leaf_307_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[22\]\[12\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xinput26 la_data_in[17] net26 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_183_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput37 la_data_in[28] net37 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_89_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_7_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_155_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10527_ _05233_ _01187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_122_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10458_ soc.cpu.PC.in\[3\] _05172_ _05173_ _05182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_237_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_217_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_48_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10389_ _05136_ _01146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_83_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12128_ _01156_ clknet_leaf_48_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[6\]\[20\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_46_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_61_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12059_ _01102_ clknet_leaf_99_wb_clk_i soc.rom_encoder_0.toggled_sram_sck vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_96_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_237_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_226_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_211_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06620_ _02356_ _02357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_168_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_80_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_244_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06551_ _02316_ _02317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_185_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_179_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05502_ soc.spi_video_ram_1.state_sram_clk_counter\[3\] _01415_ _01388_ _01416_ _01417_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_09270_ _04383_ _00779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06482_ _02214_ _02276_ _02277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_209_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08221_ soc.ram_encoder_0.output_buffer\[7\] _02563_ _03787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_147_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08152_ _03741_ _00303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_146_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_147_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07103_ _02678_ _02759_ _02760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_140_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08083_ soc.spi_video_ram_1.write_fifo.fifo_mem\[11\]\[19\] _02341_ _03691_ _03701_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_162_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07034_ _02598_ _02693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_162_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_192_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xclkbuf_leaf_195_wb_clk_i clknet_5_25_0_wb_clk_i clknet_leaf_195_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_6309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_124_wb_clk_i clknet_5_13_0_wb_clk_i clknet_leaf_124_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_103_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_216_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_130_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08985_ soc.spi_video_ram_1.write_fifo.fifo_mem\[21\]\[4\] _02399_ _04210_ _04215_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_69_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4907 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4918 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07936_ soc.spi_video_ram_1.write_fifo.fifo_mem\[12\]\[20\] soc.spi_video_ram_1.write_fifo.fifo_mem\[13\]\[20\]
+ soc.spi_video_ram_1.write_fifo.fifo_mem\[14\]\[20\] soc.spi_video_ram_1.write_fifo.fifo_mem\[15\]\[20\]
+ _02713_ _02714_ _03578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_102_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4929 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_216_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07867_ soc.spi_video_ram_1.write_fifo.fifo_mem\[15\]\[22\] _03511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09606_ soc.rom_encoder_0.input_buffer\[5\] _04584_ _04601_ _04606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06818_ _01379_ soc.ram_encoder_0.toggled_sram_sck _02489_ _02493_ _02494_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_243_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_232_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07798_ soc.spi_video_ram_1.write_fifo.fifo_mem\[29\]\[23\] _03443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_37_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09537_ _04555_ _04557_ _00873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06749_ _02430_ _00212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_71_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_227_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_212_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_244_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09468_ soc.rom_encoder_0.output_buffer\[15\] _02463_ _02464_ soc.rom_encoder_0.request_data_out\[11\]
+ _04513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_12_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_164_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_145_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_196_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08419_ soc.spi_video_ram_1.write_fifo.fifo_mem\[27\]\[7\] _02405_ _03899_ _03907_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_8_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09399_ _04458_ _00834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_36_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11430_ _00496_ clknet_leaf_37_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[30\]\[11\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_165_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_240_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_11361_ _00427_ clknet_leaf_188_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[28\]\[0\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_14_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_192_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10312_ soc.rom_loader.current_address\[10\] _05090_ _05092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_11292_ _00358_ clknet_leaf_77_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[1\]\[18\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_106_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10243_ _02250_ soc.spi_video_ram_1.write_fifo.fifo_mem\[5\]\[16\] _05041_ _05050_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_140_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_234_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_161_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_26_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_191_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10174_ _04683_ _04999_ _05006_ _03714_ _01061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_117_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_239_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_156_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_219_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_208_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_235_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_245_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_50_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_231_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_1488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11628_ _00006_ clknet_leaf_62_wb_clk_i soc.spi_video_ram_1.current_state\[1\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_128_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_1546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11559_ _00625_ clknet_leaf_298_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[25\]\[24\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_6_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_174_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_217_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_1284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05982_ soc.boot_loading_offset\[2\] _01865_ _01874_ _01875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_08770_ soc.spi_video_ram_1.write_fifo.fifo_mem\[24\]\[21\] _04061_ _04075_ _04099_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_84_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07721_ _03362_ _03363_ _03366_ _02908_ _02569_ _03367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_66_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_66_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07652_ _02902_ _03297_ _03298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_38_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_225_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_214_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06603_ _02346_ _00150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_20_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07583_ _02656_ _03220_ _03229_ _03230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_20_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06534_ _02169_ soc.spi_video_ram_1.write_fifo.fifo_mem\[0\]\[24\] _02278_ _02305_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_09322_ _02248_ soc.spi_video_ram_1.write_fifo.fifo_mem\[4\]\[15\] _04406_ _04412_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_181_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_224_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_221_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06465_ _02265_ _00093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09253_ _04374_ _00771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_181_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_222_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08204_ soc.rom_encoder_0.initializing_step\[4\] soc.rom_encoder_0.initializing_step\[3\]
+ _03772_ _03773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_72_1583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09184_ _01863_ _04333_ _04336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06396_ soc.spi_video_ram_1.fifo_in_data\[1\] _02219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_147_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_198_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08135_ _02113_ soc.spi_video_ram_1.write_fifo.fifo_mem\[10\]\[0\] _03732_ _03733_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_159_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_193_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_305_wb_clk_i clknet_5_1_0_wb_clk_i clknet_leaf_305_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_49_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08066_ _03692_ _00266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_159_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07017_ _02675_ _02676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_235_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6106 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6117 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6128 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6139 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_157_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_1444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_102_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4704 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4715 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08968_ _04205_ _00655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_44_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4726 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4737 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4748 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07919_ soc.spi_video_ram_1.write_fifo.fifo_mem\[24\]\[21\] soc.spi_video_ram_1.write_fifo.fifo_mem\[25\]\[21\]
+ soc.spi_video_ram_1.write_fifo.fifo_mem\[26\]\[21\] soc.spi_video_ram_1.write_fifo.fifo_mem\[27\]\[21\]
+ _02903_ _02904_ _03562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_4759 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08899_ _04168_ _00623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_84_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_217_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10930_ soc.spi_video_ram_1.write_fifo.fifo_mem\[8\]\[21\] _04061_ _05430_ _05454_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xclkbuf_leaf_92_wb_clk_i clknet_5_14_0_wb_clk_i clknet_leaf_92_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_131_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_56_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10861_ _01666_ _05222_ _05412_ _05417_ _01337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
Xclkbuf_leaf_21_wb_clk_i clknet_5_8_0_wb_clk_i clknet_leaf_21_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_246_1742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_213_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10792_ _05380_ _01305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_158_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_197_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_235_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_185_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_200_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_185_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_138_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11413_ _00479_ clknet_leaf_242_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[2\]\[23\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_193_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_197_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11344_ _00410_ clknet_leaf_0_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[27\]\[12\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_99_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_180_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_1590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_165_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11275_ _00341_ clknet_leaf_216_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[1\]\[1\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_152_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10226_ _02235_ soc.spi_video_ram_1.write_fifo.fifo_mem\[5\]\[9\] _05030_ _05040_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_84_1476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10157_ _02504_ _04993_ _04994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_62_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_136_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5950 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5961 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5972 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_212_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5983 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10088_ _04928_ _04939_ _04940_ _04941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_94_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5994 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_23_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_5_5_0_wb_clk_i clknet_4_2_0_wb_clk_i clknet_5_5_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_207_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_165_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_203_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_245_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_241_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_176_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06250_ soc.spi_video_ram_1.fifo_in_data\[4\] _02128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_223_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06181_ soc.video_generator_1.v_count\[8\] soc.video_generator_1.v_count\[1\] _02069_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_15_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_209_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_239_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09940_ soc.ram_encoder_0.input_bits_left\[3\] _04839_ _04843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_172_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09871_ _01598_ _04741_ _04789_ _04790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08822_ _02151_ soc.spi_video_ram_1.write_fifo.fifo_mem\[23\]\[15\] _04117_ _04128_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_115_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_230_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_246_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08753_ _04090_ _00555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_6_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05965_ _01855_ _01857_ _01858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_54_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07704_ _02581_ _03346_ _03349_ _03350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_39_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_72_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05896_ _01758_ _01761_ _01792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_08684_ soc.spi_video_ram_1.fifo_in_data\[13\] _04050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_96_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1908 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07635_ soc.spi_video_ram_1.output_buffer\[10\] _02882_ _03280_ _03281_ _03282_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_187_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_242_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_228_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07566_ _03208_ _03209_ _03212_ _02976_ _02929_ _03213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_179_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09305_ _02231_ soc.spi_video_ram_1.write_fifo.fifo_mem\[4\]\[7\] _04395_ _04403_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_55_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06517_ _02296_ _00114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_126_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07497_ _03135_ _03144_ _02567_ _03145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_186_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09236_ _02225_ soc.spi_video_ram_1.write_fifo.fifo_mem\[9\]\[4\] _04365_ _04366_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06448_ soc.spi_video_ram_1.fifo_in_address\[2\] _02254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_6_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09167_ soc.video_generator_1.v_count\[3\] _04323_ _04324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_135_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06379_ _02169_ soc.spi_video_ram_1.write_fifo.fifo_mem\[17\]\[24\] _02181_ _02208_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_202_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08118_ _01836_ _03719_ _03721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_119_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09098_ _04279_ _00711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_107_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_194_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_162_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_155_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08049_ _03683_ _00258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_150_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11060_ _00126_ clknet_leaf_43_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[0\]\[27\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_192_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_5202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_133_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_27_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10011_ soc.ram_encoder_0.request_data_out\[8\] soc.ram_encoder_0.data_out\[8\] _04889_
+ _04891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_62_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_5235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_118_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3800 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_185_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3811 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3822 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3833 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11962_ _01021_ clknet_leaf_162_wb_clk_i soc.ram_encoder_0.request_data_out\[15\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_4589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3844 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_245_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3855 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_244_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3866 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3877 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10913_ _05445_ _01361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3888 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3899 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11893_ _00952_ clknet_leaf_74_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[3\]\[19\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_60_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_232_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10844_ soc.spi_video_ram_1.fifo_in_address\[10\] _05393_ _05408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_73_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_298_wb_clk_i clknet_5_1_0_wb_clk_i clknet_leaf_298_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_13_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10775_ _04065_ _05359_ _05371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_158_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_227_wb_clk_i clknet_5_20_0_wb_clk_i clknet_leaf_227_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_201_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_158_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_220_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_205_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_173_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_157_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_126_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_181_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11327_ _00393_ clknet_leaf_298_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[26\]\[24\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_99_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_218_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11258_ _00324_ clknet_leaf_99_wb_clk_i net64 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_84_1284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10209_ _05031_ _01071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_95_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11189_ _00255_ clknet_leaf_60_wb_clk_i soc.spi_video_ram_1.output_buffer\[1\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_6481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_171_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_132_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5780 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_95_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_236_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5791 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05750_ _01556_ _01654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_54_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05681_ _01556_ _01587_ _01588_ _01589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
XFILLER_235_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_224_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07420_ _02784_ soc.spi_video_ram_1.write_fifo.fifo_mem\[10\]\[27\] _03069_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_50_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07351_ _02703_ soc.spi_video_ram_1.write_fifo.fifo_mem\[20\]\[28\] _03000_ _03001_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_182_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06302_ soc.spi_video_ram_1.fifo_in_address\[5\] _02163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_07282_ _02931_ soc.spi_video_ram_1.write_fifo.fifo_mem\[13\]\[10\] _02932_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_149_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_206_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06233_ soc.spi_video_ram_1.write_fifo.write_pointer\[4\] _02115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_09021_ _04234_ _00679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_121_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06164_ _02055_ _02056_ _02057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_85_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_06095_ _01987_ _01988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_116_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_236_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_160_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09923_ soc.rom_encoder_0.initializing_step\[3\] _04825_ soc.rom_encoder_0.initializing_step\[4\]
+ _04829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_193_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_63_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09854_ _01705_ _04740_ _04776_ _04777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_100_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08805_ _02134_ soc.spi_video_ram_1.write_fifo.fifo_mem\[23\]\[7\] _04117_ _04119_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09785_ _04722_ _00956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06997_ _02638_ _02641_ _02649_ _02654_ _02656_ _02657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XTAP_3107 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3118 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3129 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08736_ _04081_ _00547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05948_ _01836_ soc.video_generator_1.h_count\[7\] soc.video_generator_1.h_count\[6\]
+ _01840_ _01841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_67_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_226_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1705 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08667_ _04039_ _00520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_96_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05879_ _01771_ _01774_ _01776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_53_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1716 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1727 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_214_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07618_ _02704_ soc.spi_video_ram_1.write_fifo.fifo_mem\[11\]\[25\] _02593_ _03265_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1749 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08598_ _04003_ _00487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_74_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_241_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_198_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07549_ _03194_ _03195_ _02976_ _03196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_70_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_320_wb_clk_i clknet_5_0_0_wb_clk_i clknet_leaf_320_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_224_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10560_ _04243_ _05249_ _05250_ _01203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_128_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_210_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09219_ _04341_ _01819_ _04355_ _00756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_194_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10491_ soc.cpu.PC.REG.data\[11\] _05206_ _05207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_5_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_12230_ _01258_ clknet_leaf_310_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[29\]\[12\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_120_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12161_ _01189_ clknet_leaf_185_wb_clk_i soc.ram_encoder_0.address\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_100_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_135_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11112_ _00178_ clknet_leaf_285_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[12\]\[21\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_151_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12092_ _01120_ net86 soc.cpu.ALU.x\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_81_1413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_235_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5010 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11043_ _00109_ clknet_leaf_18_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[0\]\[10\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_122_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5021 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5032 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_49_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5043 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_172_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5054 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5065 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5076 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5087 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_218_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5098 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_79_1320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_4375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11945_ _01004_ clknet_leaf_161_wb_clk_i soc.ram_encoder_0.input_buffer\[11\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_166_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_217_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_206_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2940 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2951 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3696 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2962 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_127_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_233_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2973 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11876_ _00935_ clknet_leaf_258_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[3\]\[2\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2984 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2995 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_127_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_246_1391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10827_ _05399_ _01321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_242_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_203_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10758_ _03297_ _05358_ _05362_ _01289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_9_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_146_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_200_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_186_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_51_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10689_ _05309_ _05325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_103_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_142_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_206_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06920_ _00002_ _02581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_190_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_116_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_214_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06851_ soc.rom_encoder_0.output_bits_left\[3\] _02513_ _02523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_95_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05802_ _01670_ soc.cpu.ALU.x\[7\] _01703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_95_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09570_ soc.rom_encoder_0.input_bits_left\[2\] _04575_ soc.rom_encoder_0.input_bits_left\[3\]
+ _04581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_49_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06782_ _02458_ _02460_ _02461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_208_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08521_ _03961_ _00452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_82_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05733_ soc.ram_data_out\[3\] _01579_ _01638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_188_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_149_wb_clk_i clknet_5_29_0_wb_clk_i clknet_leaf_149_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_51_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08452_ soc.spi_video_ram_1.write_fifo.fifo_mem\[27\]\[23\] _02264_ _03898_ _03924_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_05664_ _01568_ _01569_ _01570_ _01571_ _01572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_145_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07403_ _03048_ _03049_ _03050_ _03051_ _02929_ _03052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_223_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08383_ _03887_ _00388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05595_ _01492_ _01503_ _01504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_177_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_220_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07334_ _02900_ _02984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_225_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_177_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07265_ _02915_ _00242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_176_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09004_ _04047_ _04225_ _04226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_118_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06216_ _01502_ _01503_ _01492_ _02102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_07196_ soc.spi_video_ram_1.write_fifo.fifo_mem\[28\]\[7\] soc.spi_video_ram_1.write_fifo.fifo_mem\[29\]\[7\]
+ soc.spi_video_ram_1.write_fifo.fifo_mem\[30\]\[7\] soc.spi_video_ram_1.write_fifo.fifo_mem\[31\]\[7\]
+ _02769_ _02770_ _02849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_219_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_192_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06147_ _01870_ _02036_ _02039_ _01847_ _02040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_145_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06078_ _01926_ _01902_ _01967_ _01970_ _01971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_116_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09906_ _04254_ _04734_ _04816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_28_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_59_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_150_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_232_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09837_ _04583_ _04761_ _04762_ _04763_ _04764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_63_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_8_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_230_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09768_ _02248_ soc.spi_video_ram_1.write_fifo.fifo_mem\[3\]\[15\] _04708_ _04714_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_100_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_185_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_227_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08719_ _03169_ _04046_ _04071_ _00540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_167_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09699_ soc.cpu.PC.REG.data\[11\] soc.rom_loader.current_address\[11\] _04638_ _04668_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_2236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_148_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11730_ _00791_ clknet_leaf_262_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[4\]\[3\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_215_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_14_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_186_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11661_ _00722_ clknet_leaf_65_wb_clk_i soc.spi_video_ram_1.state_counter\[0\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_199_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_148_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_243_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10612_ soc.spi_video_ram_1.write_fifo.fifo_mem\[19\]\[5\] _02401_ _05278_ _05284_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_11592_ _00658_ clknet_leaf_276_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[22\]\[28\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_10_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_211_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10543_ _05241_ _01195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_128_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_183_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10474_ soc.cpu.PC.REG.data\[7\] _05193_ _05194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_100_1535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_12213_ _01241_ clknet_leaf_305_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[19\]\[24\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_108_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_1171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_155_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12144_ _01172_ net88 soc.cpu.PC.REG.data\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_124_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_110_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_12075_ _01118_ clknet_leaf_99_wb_clk_i soc.rom_loader.wait_fall_clk vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_123_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11026_ _00092_ clknet_leaf_266_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[16\]\[22\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_215_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4150 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4161 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4172 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4183 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_242_wb_clk_i clknet_5_16_0_wb_clk_i clknet_leaf_242_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_75_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_209_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_185_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11928_ _00987_ clknet_leaf_85_wb_clk_i soc.rom_encoder_0.initializing_step\[3\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_75_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2770 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2781 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_205_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_146_1749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2792 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11859_ _00918_ clknet_leaf_106_wb_clk_i soc.rom_encoder_0.request_address\[4\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_162_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_202_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_1413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_192_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_201_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07050_ _02583_ _02692_ _02708_ _02602_ _02709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_12_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_220_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06001_ soc.boot_loading_offset\[0\] _01870_ _01868_ _01894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_133_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_233_1722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07952_ _03587_ _03589_ _03591_ _03593_ _02568_ _03594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_151_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06903_ soc.ram_encoder_0.request_address\[0\] _02506_ _02565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_07883_ soc.spi_video_ram_1.write_fifo.fifo_mem\[0\]\[21\] soc.spi_video_ram_1.write_fifo.fifo_mem\[1\]\[21\]
+ soc.spi_video_ram_1.write_fifo.fifo_mem\[2\]\[21\] soc.spi_video_ram_1.write_fifo.fifo_mem\[3\]\[21\]
+ _02763_ _02827_ _03526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_9_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09622_ soc.rom_encoder_0.request_write _04618_ _04619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06834_ soc.ram_encoder_0.output_bits_left\[3\] _02494_ _02509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_99_1559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_231_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_228_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_209_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09553_ _02433_ _02442_ _04565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_23_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06765_ _02434_ _02435_ _02444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_83_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_184_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08504_ _02155_ soc.spi_video_ram_1.write_fifo.fifo_mem\[28\]\[17\] _03945_ _03953_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_149_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05716_ soc.gpio_i_stored\[2\] soc.cpu.AReg.data\[0\] _01603_ _01576_ _01622_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_52_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09484_ _04520_ _04524_ _04526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06696_ soc.spi_video_ram_1.write_fifo.fifo_mem\[14\]\[4\] _02399_ _02391_ _02400_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_211_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08435_ _03915_ _00412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05647_ _01552_ soc.cpu.instruction\[5\] _01555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_12_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08366_ soc.spi_video_ram_1.write_fifo.fifo_mem\[26\]\[11\] _02414_ _03877_ _03879_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_05578_ _01472_ _01487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_07317_ _02952_ _02961_ _02966_ _02585_ _02967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_71_1478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08297_ _02138_ soc.spi_video_ram_1.write_fifo.fifo_mem\[1\]\[9\] _03831_ _03841_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_137_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07248_ _02767_ _02898_ _02831_ _02899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_125_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_191_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_46_wb_clk_i clknet_5_3_0_wb_clk_i clknet_leaf_46_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_180_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_69_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07179_ _02824_ _02826_ _02829_ _02832_ _02567_ _02833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_191_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10190_ soc.hack_clock_0.counter\[1\] soc.hack_clock_0.counter\[0\] _05019_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_117_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_246_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_189_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_74_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_169_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_46_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2000 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2011 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2022 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_210_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2033 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2044 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2055 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2066 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2077 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2088 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11713_ _00774_ clknet_leaf_9_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[9\]\[15\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_188_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2099 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_242_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_187_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_204_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11644_ _00705_ clknet_leaf_308_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[20\]\[12\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_230_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_141_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_35_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput16 io_in[32] net16 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_11575_ _00641_ clknet_leaf_34_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[22\]\[11\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_196_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xinput27 la_data_in[18] net27 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_156_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput38 la_data_in[2] net38 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_6_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10526_ soc.ram_encoder_0.address\[4\] soc.cpu.AReg.data\[4\] _05228_ _05233_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_239_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_156_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10457_ soc.cpu.PC.REG.data\[3\] _05180_ _05181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_136_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_217_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_100_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_139_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10388_ _02237_ soc.spi_video_ram_1.write_fifo.fifo_mem\[6\]\[10\] _05135_ _05136_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_97_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12127_ _01155_ clknet_leaf_74_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[6\]\[19\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_111_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12058_ net36 clknet_leaf_315_wb_clk_i soc.rom_encoder_0.data_out\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_77_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11009_ _00075_ clknet_leaf_217_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[16\]\[5\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_238_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06550_ _02315_ _02316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_240_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_234_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05501_ _01387_ soc.spi_video_ram_1.state_sram_clk_counter\[1\] soc.spi_video_ram_1.state_sram_clk_counter\[0\]
+ _01416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_33_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06481_ soc.spi_video_ram_1.write_fifo.write_pointer\[4\] _01403_ _02116_ _02276_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_60_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08220_ soc.ram_encoder_0.request_address\[6\] _02506_ _03781_ soc.ram_encoder_0.output_buffer\[3\]
+ _03786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_21_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_226_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_193_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08151_ _02136_ soc.spi_video_ram_1.write_fifo.fifo_mem\[10\]\[8\] _03732_ _03741_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_140_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07102_ soc.spi_video_ram_1.write_fifo.fifo_mem\[16\]\[3\] soc.spi_video_ram_1.write_fifo.fifo_mem\[17\]\[3\]
+ soc.spi_video_ram_1.write_fifo.fifo_mem\[18\]\[3\] soc.spi_video_ram_1.write_fifo.fifo_mem\[19\]\[3\]
+ _02681_ _02758_ _02759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_08082_ _03700_ _00274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_107_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07033_ soc.spi_video_ram_1.write_fifo.fifo_mem\[0\]\[2\] soc.spi_video_ram_1.write_fifo.fifo_mem\[1\]\[2\]
+ soc.spi_video_ram_1.write_fifo.fifo_mem\[2\]\[2\] soc.spi_video_ram_1.write_fifo.fifo_mem\[3\]\[2\]
+ _02689_ _02691_ _02692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_175_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08984_ _04214_ _00662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_192_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4908 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07935_ _02596_ _03577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_4919 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_164_wb_clk_i clknet_5_27_0_wb_clk_i clknet_leaf_164_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_99_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_244_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07866_ _02704_ soc.spi_video_ram_1.write_fifo.fifo_mem\[13\]\[22\] _03509_ _02742_
+ _03510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_84_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_186_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09605_ soc.rom_encoder_0.input_buffer\[9\] _04605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_28_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06817_ _02490_ _02492_ _02493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_56_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07797_ _02575_ soc.spi_video_ram_1.write_fifo.fifo_mem\[30\]\[23\] _03441_ _02904_
+ _03442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_77_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09536_ soc.spi_video_ram_1.write_fifo.write_pointer\[1\] _04556_ _04254_ _04557_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06748_ soc.spi_video_ram_1.write_fifo.fifo_mem\[14\]\[26\] _02270_ _02390_ _02430_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_58_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_197_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_224_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09467_ _02542_ _04511_ _04512_ _00848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06679_ _02387_ _00185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_58_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_223_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_184_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_244_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_08418_ _03906_ _00404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_145_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_205_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09398_ net12 soc.spi_video_ram_1.read_value\[3\] _04454_ _04458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_212_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08349_ soc.spi_video_ram_1.write_fifo.fifo_mem\[26\]\[3\] _02397_ _03866_ _03870_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_197_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11360_ _00426_ clknet_leaf_298_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[27\]\[28\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_138_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_1406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10311_ soc.rom_loader.current_address\[10\] _05090_ _05091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_165_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11291_ _00357_ clknet_leaf_78_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[1\]\[17\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_106_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10242_ _03419_ _05044_ _05049_ _01086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_65_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10173_ soc.ram_encoder_0.initializing_step\[2\] _05003_ _05004_ _05005_ _05006_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_82_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_232_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_234_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_222_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_216_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_182_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_1440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_8_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_223_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11627_ _00005_ clknet_leaf_62_wb_clk_i soc.spi_video_ram_1.current_state\[0\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_7_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_200_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11558_ _00624_ clknet_leaf_233_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[25\]\[23\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_144_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10509_ _05220_ _05221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_156_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11489_ _00555_ clknet_leaf_319_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[24\]\[12\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_48_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_139_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_135_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05981_ _01869_ _01873_ _01874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_26_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_214_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07720_ _02919_ soc.spi_video_ram_1.write_fifo.fifo_mem\[8\]\[24\] _03365_ _03366_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_230_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_226_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_211_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_239_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_187_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07651_ soc.spi_video_ram_1.write_fifo.fifo_mem\[31\]\[14\] _03297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xclkbuf_0_wb_clk_i wb_clk_i clknet_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_19_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06602_ soc.spi_video_ram_1.write_fifo.fifo_mem\[13\]\[22\] _02262_ _02316_ _02346_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_92_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07582_ _02707_ _03221_ _03228_ _02910_ _03229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_59_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_241_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09321_ _04411_ _00802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06533_ _02304_ _00122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_1279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_55_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_206_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_209_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_61_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_33_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09252_ _02242_ soc.spi_video_ram_1.write_fifo.fifo_mem\[9\]\[12\] _04365_ _04374_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_90_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06464_ soc.spi_video_ram_1.write_fifo.fifo_mem\[16\]\[23\] _02264_ _02216_ _02265_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_22_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_181_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08203_ soc.rom_encoder_0.initializing_step\[1\] _02459_ soc.rom_encoder_0.initializing_step\[2\]
+ _03772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09183_ soc.video_generator_1.v_count\[8\] _04334_ _04335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_72_1595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06395_ _02218_ _00070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_124_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08134_ _03731_ _03732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_88_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_198_1753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08065_ soc.spi_video_ram_1.write_fifo.fifo_mem\[11\]\[10\] _02411_ _03691_ _03692_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_88_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07016_ _02672_ _02674_ _02675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_150_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_6107 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_88_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6118 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_216_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_1314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6129 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_130_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08967_ soc.spi_video_ram_1.write_fifo.fifo_mem\[22\]\[25\] _04069_ _04177_ _04205_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_4705 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4716 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_245_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4727 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4738 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07918_ _02719_ _03560_ _03561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_5_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_187_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4749 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08898_ soc.spi_video_ram_1.write_fifo.fifo_mem\[25\]\[22\] _04063_ _04143_ _04168_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_57_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_216_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07849_ _02752_ soc.spi_video_ram_1.write_fifo.fifo_mem\[30\]\[22\] _03492_ _02895_
+ _03493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_84_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_232_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10860_ soc.ram_encoder_0.data_out\[4\] _05417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_204_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_227_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09519_ _04544_ _00868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_231_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10791_ _02219_ soc.spi_video_ram_1.write_fifo.fifo_mem\[7\]\[1\] _05378_ _05380_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_71_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_207_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_164_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_73_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_1438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xclkbuf_leaf_61_wb_clk_i clknet_5_9_0_wb_clk_i clknet_leaf_61_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XPHY_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_142_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_51_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_228_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_184_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11412_ _00478_ clknet_leaf_253_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[2\]\[22\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_240_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_201_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11343_ _00409_ clknet_leaf_34_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[27\]\[11\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_193_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_1471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11274_ _00340_ clknet_leaf_221_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[1\]\[0\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_84_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_234_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_175_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10225_ _05039_ _01079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_239_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10156_ _03778_ _04876_ _04925_ _04992_ _04993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_79_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_5940 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_5951 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5962 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_23_1726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_208_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5973 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10087_ net3 _04834_ _04940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_43_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5984 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5995 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_235_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_223_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_188_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10989_ _00055_ clknet_leaf_4_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[17\]\[14\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_43_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_206_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06180_ _02031_ _01839_ _02067_ _02068_ net75 vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_184_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_217_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09870_ _04603_ _04761_ _04762_ _04788_ _04789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_119_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_154_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08821_ _04127_ _00586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_135_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08752_ soc.spi_video_ram_1.write_fifo.fifo_mem\[24\]\[12\] _04047_ _04087_ _04090_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_227_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05964_ soc.video_generator_1.v_count\[4\] _01856_ _01857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_26_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07703_ _02590_ soc.spi_video_ram_1.write_fifo.fifo_mem\[28\]\[24\] _03348_ _02740_
+ _03349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_2_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08683_ _03140_ _04046_ _04049_ _00526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_54_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_230_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05895_ _01732_ _01733_ _01790_ _01791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_214_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_148_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07634_ _02034_ _01897_ _02625_ _02734_ _03281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_246_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1909 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_213_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07565_ _02744_ soc.spi_video_ram_1.write_fifo.fifo_mem\[8\]\[13\] _03211_ _03212_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_59_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_224_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09304_ _04402_ _00794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_94_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06516_ _02151_ soc.spi_video_ram_1.write_fifo.fifo_mem\[0\]\[15\] _02290_ _02296_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_22_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_210_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07496_ _02952_ _03136_ _03143_ _02585_ _03144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_55_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09235_ _04359_ _04365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_194_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_181_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06447_ _02253_ _00087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_22_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09166_ _04317_ _04322_ _04323_ _00735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_06378_ _02207_ _00064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_108_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08117_ _03713_ _03719_ _03720_ _00289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_135_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09097_ _02254_ soc.spi_video_ram_1.write_fifo.fifo_mem\[20\]\[18\] _04270_ _04279_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_190_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08048_ soc.spi_video_ram_1.write_fifo.fifo_mem\[11\]\[2\] _02395_ _03680_ _03683_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_235_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_172_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10010_ _04890_ _01013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_131_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09999_ _04884_ _01008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_5247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3801 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_217_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3812 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3823 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11961_ _01020_ clknet_leaf_114_wb_clk_i soc.ram_encoder_0.request_data_out\[14\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_4568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3834 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_178_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3845 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3856 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_56_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_233_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3867 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10912_ soc.spi_video_ram_1.write_fifo.fifo_mem\[8\]\[12\] _04047_ _05442_ _05445_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_3878 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11892_ _00951_ clknet_leaf_77_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[3\]\[18\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_205_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3889 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10843_ _03259_ _05392_ _05407_ _01329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_60_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_207_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_197_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10774_ _03491_ _05358_ _05370_ _01297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_13_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_200_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_164_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_185_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_220_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_267_wb_clk_i clknet_5_7_0_wb_clk_i clknet_leaf_267_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_197_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11326_ _00392_ clknet_leaf_233_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[26\]\[23\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_99_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_180_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_181_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_141_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11257_ _00323_ clknet_leaf_282_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[10\]\[28\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_49_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_214_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_171_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10208_ _02213_ soc.spi_video_ram_1.write_fifo.fifo_mem\[5\]\[0\] _05030_ _05031_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_68_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_84_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11188_ _00254_ clknet_leaf_60_wb_clk_i soc.spi_video_ram_1.output_buffer\[2\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_6471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_136_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10139_ soc.ram_encoder_0.request_data_out\[14\] _04929_ _04980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_212_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_209_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5770 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5781 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5792 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_48_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05680_ _01560_ _01584_ _01588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_165_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_149_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_225_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07350_ _02679_ soc.spi_video_ram_1.write_fifo.fifo_mem\[21\]\[28\] _03000_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_93_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_147_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06301_ _02162_ _00032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_108_1466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07281_ _02573_ _02931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_148_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09020_ soc.spi_video_ram_1.write_fifo.fifo_mem\[21\]\[20\] _02343_ _04221_ _04234_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_34_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06232_ _01400_ _01405_ _02114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_145_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06163_ _01849_ _01939_ _02034_ _01940_ _02056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_89_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06094_ _01902_ _01969_ _01987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_85_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_171_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09922_ _04243_ _04826_ _04828_ _00987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_176_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09853_ _04594_ _04761_ _04762_ _04775_ _04776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_8_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08804_ _04118_ _00578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_100_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_246_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09784_ _02264_ soc.spi_video_ram_1.write_fifo.fifo_mem\[3\]\[23\] _04696_ _04722_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_100_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06996_ _02655_ _02656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_3108 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3119 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08735_ soc.spi_video_ram_1.write_fifo.fifo_mem\[24\]\[4\] _02399_ _04076_ _04081_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_05947_ _01838_ _01839_ _01840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_100_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_215_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08666_ soc.spi_video_ram_1.write_fifo.fifo_mem\[15\]\[6\] _02403_ _04032_ _04039_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_05878_ _01771_ _01774_ _01775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_22_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_187_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_242_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1717 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07617_ _03047_ soc.spi_video_ram_1.write_fifo.fifo_mem\[10\]\[25\] _03264_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_1728 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1739 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08597_ _02124_ soc.spi_video_ram_1.write_fifo.fifo_mem\[30\]\[2\] _04000_ _04003_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_179_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_5_31_0_wb_clk_i clknet_4_15_0_wb_clk_i clknet_5_31_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_07548_ _02926_ soc.spi_video_ram_1.write_fifo.fifo_mem\[16\]\[13\] _03195_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_74_1487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07479_ soc.spi_video_ram_1.write_fifo.fifo_mem\[0\]\[12\] soc.spi_video_ram_1.write_fifo.fifo_mem\[1\]\[12\]
+ soc.spi_video_ram_1.write_fifo.fifo_mem\[2\]\[12\] soc.spi_video_ram_1.write_fifo.fifo_mem\[3\]\[12\]
+ _02919_ _02577_ _03127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_50_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_167_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09218_ _04050_ _04346_ _04355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_10490_ _04664_ _05203_ _05206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_108_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_202_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09149_ _04294_ _04310_ _00731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_159_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_146_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12160_ _01188_ clknet_leaf_149_wb_clk_i soc.ram_encoder_0.address\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_194_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_162_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_155_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11111_ _00177_ clknet_leaf_50_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[12\]\[20\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_85_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12091_ soc.cpu.PC.in\[14\] net89 soc.cpu.AReg.data\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_150_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5000 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11042_ _00108_ clknet_leaf_247_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[0\]\[9\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_5011 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5022 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_231_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5033 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5044 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5055 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5066 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_213_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_4332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5077 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5088 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5099 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11944_ _01003_ clknet_leaf_160_wb_clk_i soc.ram_encoder_0.input_buffer\[10\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2930 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2941 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2952 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3697 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2963 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_232_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_229_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11875_ _00934_ clknet_leaf_215_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[3\]\[1\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2974 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2985 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2996 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10826_ _02252_ soc.spi_video_ram_1.write_fifo.fifo_mem\[7\]\[17\] _05389_ _05399_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_60_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_186_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_201_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_158_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10757_ _04052_ _05359_ _05362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_125_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_105_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_187_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_220_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10688_ _05321_ _05324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_139_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_173_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_153_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11309_ _00375_ clknet_leaf_201_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[26\]\[6\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_218_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12289_ _01317_ clknet_leaf_312_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[7\]\[13\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_136_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06850_ _02445_ _02515_ _02520_ _02521_ _02522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_68_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_228_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05801_ _01557_ _01702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_83_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06781_ _02459_ _02449_ _02460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_222_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08520_ _02171_ soc.spi_video_ram_1.write_fifo.fifo_mem\[28\]\[25\] _03933_ _03961_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_05732_ _01557_ _01636_ _01637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_36_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_224_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08451_ _03923_ _00420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05663_ soc.cpu.AReg.data\[9\] soc.cpu.AReg.data\[8\] _01571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_184_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07402_ _02922_ soc.spi_video_ram_1.write_fifo.fifo_mem\[9\]\[11\] _03024_ _03051_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08382_ soc.spi_video_ram_1.write_fifo.fifo_mem\[26\]\[19\] _02341_ _03877_ _03887_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_162_1722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05594_ _01501_ soc.spi_video_ram_1.output_buffer\[22\] _01477_ soc.spi_video_ram_1.output_buffer\[23\]
+ _01503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_182_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_189_wb_clk_i clknet_5_22_0_wb_clk_i clknet_leaf_189_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_36_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07333_ _02970_ _02977_ _02982_ _02983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_91_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_177_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_118_wb_clk_i clknet_5_26_0_wb_clk_i clknet_leaf_118_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_137_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07264_ soc.spi_video_ram_1.output_buffer\[14\] _02914_ _02633_ _02915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_137_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09003_ _04209_ _04225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_06215_ _02091_ _02098_ _02099_ _02100_ _02101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_178_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07195_ _01507_ _02676_ _02845_ _02848_ _00239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_118_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06146_ _01949_ _01893_ _02037_ _02038_ _02039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or4_1
XFILLER_30_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06077_ _01891_ _01969_ _01970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_132_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09905_ _02443_ _04809_ _04815_ _04254_ _00983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_160_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09836_ soc.rom_encoder_0.request_data_out\[4\] _04743_ _04763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_101_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_150_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_210_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09767_ _04713_ _00947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_73_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06979_ soc.spi_video_ram_1.write_fifo.fifo_mem\[12\]\[1\] soc.spi_video_ram_1.write_fifo.fifo_mem\[13\]\[1\]
+ soc.spi_video_ram_1.write_fifo.fifo_mem\[14\]\[1\] soc.spi_video_ram_1.write_fifo.fifo_mem\[15\]\[1\]
+ _02607_ _02636_ _02639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_74_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08718_ _03927_ _04048_ _04071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09698_ _04618_ _04666_ _04667_ _00924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_2226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08649_ _04029_ _00512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_70_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_214_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_148_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11660_ _00721_ clknet_leaf_276_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[20\]\[28\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_35_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_230_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_70_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_208_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_70_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10611_ _05283_ _01221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_126_1352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11591_ _00657_ clknet_leaf_44_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[22\]\[27\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_70_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_210_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10542_ soc.ram_encoder_0.address\[12\] soc.cpu.AReg.data\[12\] _05227_ _05241_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_161_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_194_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_210_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10473_ soc.cpu.PC.REG.data\[5\] soc.cpu.PC.REG.data\[6\] _05186_ _05193_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_68_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12212_ _01240_ clknet_leaf_234_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[19\]\[23\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_124_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12143_ _01171_ net88 soc.cpu.PC.REG.data\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_124_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_235_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12074_ _01117_ clknet_leaf_110_wb_clk_i soc.rom_loader.current_address\[14\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_96_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11025_ _00091_ clknet_leaf_236_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[16\]\[21\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_46_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_77_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4140 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_237_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_150_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4151 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_4162 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_111_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4173 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4184 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_206_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11927_ _00986_ clknet_leaf_86_wb_clk_i soc.rom_encoder_0.initializing_step\[2\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_79_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_233_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2760 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2771 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2782 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_127_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_226_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2793 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_127_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11858_ _00917_ clknet_leaf_108_wb_clk_i soc.rom_encoder_0.request_address\[3\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_242_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xclkbuf_leaf_282_wb_clk_i clknet_5_7_0_wb_clk_i clknet_leaf_282_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_183_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10809_ _05377_ _05389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_159_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11789_ _00850_ clknet_leaf_63_wb_clk_i soc.spi_video_ram_1.buffer_index\[0\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_14_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_211_wb_clk_i clknet_5_20_0_wb_clk_i clknet_leaf_211_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_174_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06000_ soc.video_generator_1.h_count\[4\] _01891_ _01892_ _01893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_127_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_31_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_154_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_86_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07951_ _02571_ _03592_ _02602_ _03593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_114_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_190_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06902_ _02556_ _02562_ _02564_ _00231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07882_ _03525_ _00249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_229_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_214_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_1505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_233_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06833_ _02500_ _02497_ _02506_ _02507_ _02508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
X_09621_ _04617_ _04618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_95_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09552_ _04564_ _00881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06764_ _02433_ _02442_ _02443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_24_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08503_ _03952_ _00443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_149_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05715_ net79 _01564_ _01576_ _01577_ _01621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_37_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09483_ _01518_ _04520_ _04524_ _04525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_52_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06695_ soc.spi_video_ram_1.fifo_in_data\[4\] _02399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_145_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08434_ soc.spi_video_ram_1.write_fifo.fifo_mem\[27\]\[14\] _02246_ _03910_ _03915_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_51_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05646_ soc.cpu.DMuxJMP.sel\[0\] _01554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_93_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_212_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_180_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08365_ _03878_ _00379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05577_ _01462_ _01485_ _01486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_225_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_240_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_211_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07316_ _02962_ _02963_ _02965_ _02722_ _02900_ _02966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_108_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_20_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08296_ _03840_ _00348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_176_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07247_ soc.spi_video_ram_1.write_fifo.fifo_mem\[24\]\[9\] soc.spi_video_ram_1.write_fifo.fifo_mem\[25\]\[9\]
+ soc.spi_video_ram_1.write_fifo.fifo_mem\[26\]\[9\] soc.spi_video_ram_1.write_fifo.fifo_mem\[27\]\[9\]
+ _02893_ _02827_ _02898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_192_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_164_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07178_ _02650_ _02830_ _02831_ _02832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_145_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_238_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06129_ _01967_ _01922_ _02021_ _02022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_106_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_86_wb_clk_i clknet_5_14_0_wb_clk_i clknet_leaf_86_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_156_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_15_wb_clk_i clknet_5_2_0_wb_clk_i clknet_leaf_15_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_28_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_232_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_219_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_169_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09819_ net6 _04566_ _04749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_100_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2001 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2012 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2023 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2034 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_160_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2045 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2056 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_215_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_188_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2067 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2078 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11712_ _00773_ clknet_leaf_7_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[9\]\[14\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2089 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_199_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_243_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11643_ _00704_ clknet_leaf_36_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[20\]\[11\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_196_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_180_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_211_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11574_ _00640_ clknet_leaf_20_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[22\]\[10\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xinput17 io_in[33] net17 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_204_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput28 la_data_in[19] net28 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_183_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput39 la_data_in[3] net39 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_10525_ _05232_ _01186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_122_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10456_ soc.cpu.PC.REG.data\[0\] soc.cpu.PC.REG.data\[1\] soc.cpu.PC.REG.data\[2\]
+ _05180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_108_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10387_ _05122_ _05135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_124_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12126_ _01154_ clknet_leaf_79_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[6\]\[18\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_35_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_12057_ net35 clknet_leaf_173_wb_clk_i soc.rom_encoder_0.data_out\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_42_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_215_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11008_ _00074_ clknet_leaf_140_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[16\]\[4\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_113_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_37_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_209_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_1435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05500_ soc.spi_video_ram_1.state_sram_clk_counter\[2\] _01415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_55_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06480_ _02275_ _00098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_61_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_33_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_18_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_187_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08150_ _03740_ _00302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_119_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_222_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_174_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07101_ _02598_ _02758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_119_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08081_ soc.spi_video_ram_1.write_fifo.fifo_mem\[11\]\[18\] _02339_ _03691_ _03700_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_105_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_220_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07032_ _02690_ _02691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_175_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_174_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_196_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xclkbuf_3_0_0_wb_clk_i clknet_2_0_0_wb_clk_i clknet_3_0_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_157_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_103_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_244_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08983_ soc.spi_video_ram_1.write_fifo.fifo_mem\[21\]\[3\] _02397_ _04210_ _04214_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_87_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_233_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07934_ _02678_ _03575_ _03576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_130_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4909 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07865_ _02907_ soc.spi_video_ram_1.write_fifo.fifo_mem\[12\]\[22\] _03509_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_111_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_228_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09604_ _04603_ _04585_ _04604_ _00893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06816_ _02480_ _02491_ _02492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_42_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07796_ _03054_ _03440_ _03441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_83_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_244_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06747_ _02429_ _00211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09535_ _01444_ _04552_ _04556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XPHY_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_184_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09466_ soc.rom_encoder_0.output_buffer\[18\] _04479_ _04512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_06678_ _02177_ soc.spi_video_ram_1.write_fifo.fifo_mem\[12\]\[28\] _02356_ _02387_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_52_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_145_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08417_ soc.spi_video_ram_1.write_fifo.fifo_mem\[27\]\[6\] _02403_ _03899_ _03906_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_106_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05629_ soc.spi_video_ram_1.buffer_index\[4\] _01529_ _01537_ _01538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_240_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09397_ _04457_ _00833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_178_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08348_ _03869_ _00371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_162_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_205_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08279_ _02113_ soc.spi_video_ram_1.write_fifo.fifo_mem\[1\]\[0\] _03831_ _03832_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_165_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10310_ _05071_ _05089_ _05090_ _01112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_180_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_193_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_165_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11290_ _00356_ clknet_leaf_77_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[1\]\[16\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_98_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10241_ soc.spi_video_ram_1.fifo_in_data\[15\] _05045_ _05049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_175_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10172_ soc.ram_encoder_0.initializing_step\[2\] soc.ram_encoder_0.initializing_step\[1\]
+ soc.ram_encoder_0.initializing_step\[0\] _05005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_136_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_160_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_152_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_82_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_21_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_210_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_234_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_187_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_179_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_230_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11626_ _00692_ clknet_leaf_32_wb_clk_i _00004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_30_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11557_ _00623_ clknet_leaf_251_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[25\]\[22\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_239_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_221_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10508_ _01455_ _05219_ _05220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_128_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11488_ _00554_ clknet_leaf_33_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[24\]\[11\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_109_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10439_ soc.cpu.DMuxJMP.sel\[1\] _05166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_87_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_174_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12109_ _01137_ clknet_leaf_245_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[6\]\[1\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_97_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05980_ soc.boot_loading_offset\[0\] _01869_ _01870_ _01872_ _01873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XTAP_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_238_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07650_ soc.spi_video_ram_1.write_fifo.fifo_mem\[24\]\[14\] soc.spi_video_ram_1.write_fifo.fifo_mem\[25\]\[14\]
+ soc.spi_video_ram_1.write_fifo.fifo_mem\[26\]\[14\] soc.spi_video_ram_1.write_fifo.fifo_mem\[27\]\[14\]
+ _02902_ _02894_ _03296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_65_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_226_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06601_ _02345_ _00149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_4_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07581_ _02582_ _03224_ _03227_ _03228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_230_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_240_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09320_ _02246_ soc.spi_video_ram_1.write_fifo.fifo_mem\[4\]\[14\] _04406_ _04411_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06532_ _02167_ soc.spi_video_ram_1.write_fifo.fifo_mem\[0\]\[23\] _02278_ _02304_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_55_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_181_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09251_ _04373_ _00770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06463_ soc.spi_video_ram_1.fifo_in_address\[7\] _02264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_222_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08202_ _03764_ _03768_ _03769_ _03770_ _03771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_09182_ _04331_ _04332_ _04334_ _04317_ _00740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_193_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_147_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06394_ soc.spi_video_ram_1.write_fifo.fifo_mem\[16\]\[0\] _02213_ _02217_ _02218_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_159_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08133_ _03730_ _03731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_105_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_162_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08064_ _03678_ _03691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_159_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_162_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07015_ net18 _02673_ _02674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_150_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_200_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_190_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_6108 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_89_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_6119 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_5407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_192_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08966_ _04204_ _00654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_103_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4706 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4717 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4728 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07917_ _02952_ _03556_ _03559_ _03560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_97_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4739 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08897_ _04167_ _00622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_56_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xclkbuf_leaf_314_wb_clk_i clknet_5_1_0_wb_clk_i clknet_leaf_314_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_229_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_17_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07848_ _03139_ _03491_ _03492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_57_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_229_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_245_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_216_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07779_ _02656_ _03414_ _03423_ _03424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_71_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_207_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09518_ _02272_ soc.cpu.AReg.data\[11\] _01459_ _04544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_10790_ _05379_ _01304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_129_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09449_ soc.rom_encoder_0.output_buffer\[15\] _04479_ _04498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_158_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_185_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_160_1319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_212_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_16_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11411_ _00477_ clknet_leaf_230_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[2\]\[21\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_71_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11342_ _00408_ clknet_leaf_17_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[27\]\[10\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_181_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_30_wb_clk_i clknet_5_9_0_wb_clk_i clknet_leaf_30_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_11273_ _00339_ clknet_leaf_168_wb_clk_i soc.ram_encoder_0.output_buffer\[19\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_181_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10224_ _02233_ soc.spi_video_ram_1.write_fifo.fifo_mem\[5\]\[8\] _05030_ _05039_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_45_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10155_ _02499_ _02551_ _04991_ _04992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XTAP_5930 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5941 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_216_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5952 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5963 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10086_ soc.ram_encoder_0.request_data_out\[2\] _04930_ _04939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_5974 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5985 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_87_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_5996 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_130_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_208_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_222_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_235_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10988_ _00054_ clknet_leaf_39_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[17\]\[13\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_200_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_204_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_182_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_188_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_198_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11609_ _00675_ clknet_leaf_26_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[21\]\[16\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_15_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_141_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_176_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_213_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08820_ _02149_ soc.spi_video_ram_1.write_fifo.fifo_mem\[23\]\[14\] _04117_ _04127_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_140_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_234_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05963_ soc.video_generator_1.v_count\[7\] _01849_ soc.video_generator_1.v_count\[5\]
+ _01856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_08751_ _04089_ _00554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_239_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_152_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07702_ _02573_ _03347_ _03348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_66_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_187_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05894_ _01787_ _01789_ _01790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_08682_ _04047_ _04048_ _04049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_93_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_241_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_227_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_246_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07633_ _03231_ _03278_ _03279_ _03280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_241_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_198_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07564_ _03139_ _03210_ _03211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_5_21_0_wb_clk_i clknet_4_10_0_wb_clk_i clknet_5_21_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_80_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06515_ _02295_ _00113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09303_ _02229_ soc.spi_video_ram_1.write_fifo.fifo_mem\[4\]\[6\] _04395_ _04402_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_110_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07495_ _03137_ _03138_ _02900_ _03142_ _03143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_55_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09234_ _04364_ _00762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06446_ soc.spi_video_ram_1.write_fifo.fifo_mem\[16\]\[17\] _02252_ _02238_ _02253_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_72_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_33_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_210_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09165_ soc.video_generator_1.v_count\[2\] _04321_ _04323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_06377_ _02167_ soc.spi_video_ram_1.write_fifo.fifo_mem\[17\]\[23\] _02181_ _02207_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_175_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_222_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08116_ soc.video_generator_1.h_count\[4\] _03717_ _03720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_135_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09096_ _04278_ _00710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_190_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08047_ _03682_ _00257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_150_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_172_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09998_ soc.ram_encoder_0.request_data_out\[2\] soc.ram_encoder_0.data_out\[2\] _04880_
+ _04884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_237_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_213_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08949_ soc.spi_video_ram_1.write_fifo.fifo_mem\[22\]\[16\] _02335_ _04189_ _04196_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_9_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3802 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3813 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11960_ _01019_ clknet_leaf_162_wb_clk_i soc.ram_encoder_0.request_data_out\[13\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_4569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3824 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3835 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3846 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3857 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10911_ _05444_ _01360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3868 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3879 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11891_ _00950_ clknet_leaf_78_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[3\]\[17\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_204_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_217_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10842_ soc.spi_video_ram_1.fifo_in_address\[9\] _05393_ _05407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_72_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_240_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_92_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10773_ _04063_ _05359_ _05370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_9_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_199_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_240_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_201_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_1488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_177_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_153_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11325_ _00391_ clknet_leaf_251_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[26\]\[22\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_181_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11256_ _00322_ clknet_leaf_271_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[10\]\[27\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_134_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_236_wb_clk_i clknet_5_5_0_wb_clk_i clknet_leaf_236_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_122_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10207_ _05029_ _05030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_68_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11187_ _00253_ clknet_leaf_58_wb_clk_i soc.spi_video_ram_1.output_buffer\[3\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_6450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10138_ _04952_ _04979_ _01051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_6494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_227_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5760 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5771 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5782 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_114_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5793 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10069_ _02503_ _04679_ _04834_ _04836_ _04924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_23_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_209_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_223_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_210_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_206_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06300_ _02161_ soc.spi_video_ram_1.write_fifo.fifo_mem\[18\]\[20\] _02119_ _02162_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_91_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07280_ _02921_ _02923_ _02925_ _02928_ _02929_ _02930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_86_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_06231_ soc.spi_video_ram_1.fifo_in_data\[0\] _02113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_117_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06162_ _01853_ soc.video_generator_1.v_count\[7\] _02055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_116_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06093_ _01891_ _01905_ _01986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_102_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09921_ _02454_ _04827_ _04818_ _04828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_217_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09852_ soc.rom_encoder_0.request_data_out\[8\] _04742_ _04775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_154_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_113_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_219_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08803_ _02132_ soc.spi_video_ram_1.write_fifo.fifo_mem\[23\]\[6\] _04117_ _04118_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_140_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09783_ _04721_ _00955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_132_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_26_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06995_ _00004_ _02655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_39_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3109 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08734_ _04080_ _00546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05946_ soc.video_generator_1.h_count\[8\] soc.video_generator_1.h_count\[9\] _01839_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_85_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_230_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05877_ _01705_ _01773_ _01774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_08665_ _04038_ _00519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_57_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1707 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_199_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07616_ _02767_ _03255_ _03262_ _02719_ _03263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_1718 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1729 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_183_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08596_ _04002_ _00486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_109_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_243_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_224_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_165_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07547_ _02920_ soc.spi_video_ram_1.write_fifo.fifo_mem\[17\]\[13\] _03194_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_243_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07478_ _03116_ _03125_ _03126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_194_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_1409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09217_ _04341_ _01803_ _04354_ _00755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06429_ _02241_ _00081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_241_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_182_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09148_ soc.spi_video_ram_1.state_counter\[9\] _04308_ _04310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_147_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09079_ _04269_ _00702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_120_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_123_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11110_ _00176_ clknet_leaf_31_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[12\]\[19\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12090_ soc.cpu.PC.in\[13\] net89 soc.cpu.AReg.data\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_172_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11041_ _00107_ clknet_leaf_220_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[0\]\[8\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_5001 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_104_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5012 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_89_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5023 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5034 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_4300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_209_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_190_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_5045 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5056 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5067 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_5078 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_5089 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_4366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_233_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11943_ _01002_ clknet_leaf_159_wb_clk_i soc.ram_encoder_0.input_buffer\[9\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_4399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2920 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2931 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_205_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2942 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2953 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3698 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11874_ _00933_ clknet_leaf_221_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[3\]\[0\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2964 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_221_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2975 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2986 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2997 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10825_ _05398_ _01320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_207_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_1743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_144_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10756_ _03199_ _05358_ _05361_ _01288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_38_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_187_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10687_ _05323_ _01257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_16_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_220_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_4_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_236_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11308_ _00374_ clknet_leaf_188_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[26\]\[5\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12288_ _01316_ clknet_leaf_308_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[7\]\[12\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_113_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_214_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11239_ _00305_ clknet_leaf_13_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[10\]\[10\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_68_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_171_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05800_ _01689_ _01694_ _01585_ _01696_ _01701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_06780_ soc.rom_encoder_0.initializing_step\[0\] _02459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_3_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_76_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05731_ _01558_ soc.cpu.ALU.x\[3\] _01636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_110_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05662_ soc.cpu.AReg.data\[14\] soc.cpu.AReg.data\[13\] _01570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_08450_ soc.spi_video_ram_1.write_fifo.fifo_mem\[27\]\[22\] _02262_ _03898_ _03923_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_91_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07401_ _02971_ soc.spi_video_ram_1.write_fifo.fifo_mem\[8\]\[11\] _03050_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_08381_ _03886_ _00387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_225_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05593_ _01501_ soc.spi_video_ram_1.output_buffer\[20\] _01477_ soc.spi_video_ram_1.output_buffer\[21\]
+ _01502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_211_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07332_ _02978_ _02979_ _02980_ _02981_ _02569_ _02982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_71_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_176_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07263_ _02058_ _02625_ _02913_ _02914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_177_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09002_ _04221_ _04224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_06214_ _01472_ _01495_ _02091_ _02100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_07194_ _01411_ _02633_ _02847_ _02848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_118_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_191_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xclkbuf_leaf_158_wb_clk_i clknet_5_27_0_wb_clk_i clknet_leaf_158_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_06145_ _01853_ soc.video_generator_1.v_count\[7\] _01959_ _02038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_121_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_160_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06076_ _01968_ _01904_ _01905_ _01969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_160_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09904_ _04812_ _04809_ soc.rom_encoder_0.current_state\[2\] _04815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_8_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09835_ _04739_ _04762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_154_1284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09766_ _02246_ soc.spi_video_ram_1.write_fifo.fifo_mem\[3\]\[14\] _04708_ _04713_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_27_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06978_ _02583_ _02637_ _02638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_08717_ _03270_ _04046_ _04070_ _00539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_2205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_215_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05929_ _01618_ soc.cpu.AReg.data\[14\] _01718_ soc.ram_data_out\[14\] _01823_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_09697_ soc.rom_encoder_0.request_address\[10\] _04618_ _04667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_242_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08648_ _02175_ soc.spi_video_ram_1.write_fifo.fifo_mem\[30\]\[27\] _03999_ _04029_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XPHY_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_203_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08579_ _03992_ _00479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_25_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_168_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10610_ soc.spi_video_ram_1.write_fifo.fifo_mem\[19\]\[4\] _02399_ _05278_ _05283_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_23_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11590_ _00656_ clknet_leaf_281_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[22\]\[26\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_204_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_195_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10541_ _05240_ _01194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_126_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_202_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10472_ _05171_ _05191_ _05192_ _01172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_178_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_139_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12211_ _01239_ clknet_leaf_252_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[19\]\[22\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_87_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_203_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_194_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_159_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_191_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_237_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12142_ _01170_ net88 soc.cpu.PC.REG.data\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_159_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12073_ _01116_ clknet_leaf_102_wb_clk_i soc.rom_loader.current_address\[13\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_85_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_215_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_151_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_238_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11024_ _00090_ clknet_leaf_263_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[16\]\[20\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_133_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4130 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4141 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4152 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4163 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4174 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4185 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_4_2_0_wb_clk_i clknet_3_1_0_wb_clk_i clknet_4_2_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_46_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11926_ _00985_ clknet_leaf_97_wb_clk_i soc.rom_encoder_0.initializing_step\[1\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XTAP_3484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2750 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_244_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2761 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2772 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2783 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11857_ _00916_ clknet_leaf_92_wb_clk_i soc.rom_encoder_0.request_address\[2\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_166_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2794 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_162_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_220_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10808_ _05388_ _01313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_158_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11788_ _00849_ clknet_leaf_101_wb_clk_i soc.rom_encoder_0.output_buffer\[19\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_53_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10739_ _05351_ _01281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_173_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xclkbuf_leaf_251_wb_clk_i clknet_5_7_0_wb_clk_i clknet_leaf_251_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_115_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_192_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07950_ soc.spi_video_ram_1.write_fifo.fifo_mem\[20\]\[20\] soc.spi_video_ram_1.write_fifo.fifo_mem\[21\]\[20\]
+ soc.spi_video_ram_1.write_fifo.fifo_mem\[22\]\[20\] soc.spi_video_ram_1.write_fifo.fifo_mem\[23\]\[20\]
+ _02769_ _02770_ _03592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_9_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_233_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06901_ soc.ram_encoder_0.output_buffer\[2\] _02563_ _02564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_96_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07881_ soc.spi_video_ram_1.output_buffer\[7\] _03524_ _02633_ _03525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_228_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09620_ _04616_ _04617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_42_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06832_ _02477_ soc.ram_encoder_0.output_bits_left\[2\] _02507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_96_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_244_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09551_ _04254_ _04255_ _04564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_06763_ soc.rom_encoder_0.current_state\[2\] _02436_ _02442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_110_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08502_ _02153_ soc.spi_video_ram_1.write_fifo.fifo_mem\[28\]\[16\] _03945_ _03952_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_224_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05714_ soc.ram_data_out\[2\] _01579_ _01563_ _01620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_36_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06694_ _02398_ _00189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09482_ _01428_ _01485_ _04524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_184_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08433_ _03914_ _00411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_58_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05645_ _01552_ _01553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_08364_ soc.spi_video_ram_1.write_fifo.fifo_mem\[26\]\[10\] _02411_ _03877_ _03878_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_05576_ _01461_ soc.spi_video_ram_1.buffer_index\[1\] _01485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_51_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07315_ _02703_ soc.spi_video_ram_1.write_fifo.fifo_mem\[28\]\[10\] _02964_ _02965_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_221_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08295_ _02136_ soc.spi_video_ram_1.write_fifo.fifo_mem\[1\]\[8\] _03831_ _03840_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_203_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07246_ _02570_ _02896_ _02897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_07177_ _02585_ _02831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_195_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06128_ _01902_ _02015_ _02020_ _02021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_65_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_219_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06059_ _01950_ _01951_ _01952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_28_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_101_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09818_ soc.rom_encoder_0.request_data_out\[1\] _04743_ _04748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_8_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_210_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_55_wb_clk_i clknet_5_24_0_wb_clk_i clknet_leaf_55_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_41_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_246_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09749_ _02229_ soc.spi_video_ram_1.write_fifo.fifo_mem\[3\]\[6\] _04697_ _04704_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_2002 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2013 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2024 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_243_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2035 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2046 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2057 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2068 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11711_ _00772_ clknet_leaf_8_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[9\]\[13\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2079 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_167_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_1317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_230_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_208_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_202_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11642_ _00703_ clknet_leaf_14_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[20\]\[10\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_14_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11573_ _00639_ clknet_leaf_254_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[22\]\[9\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_106_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput18 la_data_in[0] net18 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_128_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput29 la_data_in[1] net29 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_10524_ soc.ram_encoder_0.address\[3\] soc.cpu.AReg.data\[3\] _05228_ _05232_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_7_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xcaravel_hack_soc_220 wbs_dat_o[28] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_10455_ _05171_ _05178_ _05179_ _01168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_183_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_182_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_6_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10386_ _05134_ _01145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_174_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_151_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12125_ _01153_ clknet_leaf_80_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[6\]\[17\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_96_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12056_ net34 clknet_leaf_106_wb_clk_i soc.rom_encoder_0.data_out\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_46_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_42_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_133_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11007_ _00073_ clknet_leaf_138_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[16\]\[3\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_81_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_237_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_226_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_53_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_206_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_46_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_233_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_1447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_185_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11909_ _00968_ clknet_leaf_121_wb_clk_i soc.cpu.instruction\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_55_1409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_20_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_221_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1890 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07100_ _02710_ _02748_ _02756_ _02757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_179_1313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08080_ _03699_ _00273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_105_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_228_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_200_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07031_ _02576_ _02690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_122_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08982_ _04213_ _00661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_157_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07933_ soc.spi_video_ram_1.write_fifo.fifo_mem\[8\]\[20\] soc.spi_video_ram_1.write_fifo.fifo_mem\[9\]\[20\]
+ soc.spi_video_ram_1.write_fifo.fifo_mem\[10\]\[20\] soc.spi_video_ram_1.write_fifo.fifo_mem\[11\]\[20\]
+ _02717_ _02682_ _03575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_229_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07864_ _02643_ _03500_ _03507_ _02719_ _03508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_110_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09603_ soc.rom_encoder_0.input_buffer\[4\] _04584_ _04601_ _04604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_186_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06815_ soc.ram_encoder_0.current_state\[1\] _02491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_07795_ soc.spi_video_ram_1.write_fifo.fifo_mem\[31\]\[23\] _03440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_84_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09534_ _01441_ _04552_ _04555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_225_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06746_ soc.spi_video_ram_1.write_fifo.fifo_mem\[14\]\[25\] _02268_ _02390_ _02429_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_58_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09465_ soc.rom_encoder_0.output_buffer\[14\] _02455_ _04510_ _02461_ _04511_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_58_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_06677_ _02386_ _00184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_212_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_08416_ _03905_ _00403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05628_ _01516_ _01531_ _01533_ _01519_ _01523_ _01536_ _01537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_09396_ net11 soc.spi_video_ram_1.read_value\[2\] _04454_ _04457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_12_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_225_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_240_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_173_wb_clk_i clknet_opt_5_0_wb_clk_i clknet_leaf_173_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_71_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08347_ soc.spi_video_ram_1.write_fifo.fifo_mem\[26\]\[2\] _02395_ _03866_ _03869_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_05559_ _01467_ _01468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_193_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_102_wb_clk_i clknet_5_15_0_wb_clk_i clknet_leaf_102_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_71_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08278_ _03830_ _03831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_165_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_192_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_158_1408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_101_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07229_ _02870_ _02880_ _02626_ _02881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_49_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10240_ _03320_ _05044_ _05048_ _01085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_238_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10171_ _02485_ _05003_ _05004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_78_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_216_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_191_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_82_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_232_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_173_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_219_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_208_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_28_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_215_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_231_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_188_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_203_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_180_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_187_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11625_ _00691_ clknet_leaf_32_wb_clk_i _00003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_106_1532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_204_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_184_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11556_ _00622_ clknet_leaf_230_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[25\]\[21\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10507_ _05218_ _05015_ _05019_ _05219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_7_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11487_ _00553_ clknet_leaf_17_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[24\]\[10\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_183_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10438_ _01834_ _05164_ _01554_ _05165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_174_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10369_ _02219_ soc.spi_video_ram_1.write_fifo.fifo_mem\[6\]\[1\] _05124_ _05126_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_97_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12108_ _01136_ clknet_leaf_245_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[6\]\[0\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_112_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_215_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_230_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12039_ _01098_ clknet_leaf_273_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[5\]\[27\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_111_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_230_1749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06600_ soc.spi_video_ram_1.write_fifo.fifo_mem\[13\]\[21\] _02260_ _02316_ _02345_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_207_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07580_ _02924_ soc.spi_video_ram_1.write_fifo.fifo_mem\[4\]\[13\] _03226_ _02927_
+ _03227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_80_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_5_11_0_wb_clk_i clknet_4_5_0_wb_clk_i clknet_5_11_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_94_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_146_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06531_ _02303_ _00121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_94_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_179_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_228_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_0_wb_clk_i clknet_5_0_0_wb_clk_i clknet_leaf_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_22_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09250_ _02240_ soc.spi_video_ram_1.write_fifo.fifo_mem\[9\]\[11\] _04365_ _04373_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_94_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06462_ _02263_ _00092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_146_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08201_ soc.rom_encoder_0.output_buffer\[16\] _03770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_06393_ _02216_ _02217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_09181_ _01856_ _04333_ _04334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_222_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_187_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_239_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08132_ _02114_ _03729_ _03730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_159_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_135_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_147_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08063_ _03690_ _00265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_162_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07014_ soc.spi_video_ram_1.current_state\[0\] _01411_ _02673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_190_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_108_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_6109 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_170_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08965_ soc.spi_video_ram_1.write_fifo.fifo_mem\[22\]\[24\] _04067_ _04177_ _04204_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_233_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4707 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4718 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_170_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07916_ _02689_ soc.spi_video_ram_1.write_fifo.fifo_mem\[20\]\[21\] _03558_ _02742_
+ _03559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_4729 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_151_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08896_ soc.spi_video_ram_1.write_fifo.fifo_mem\[25\]\[21\] _04061_ _04143_ _04167_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_111_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_25_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07847_ soc.spi_video_ram_1.write_fifo.fifo_mem\[31\]\[22\] _03491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_84_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_244_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_186_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07778_ _02707_ _03415_ _03422_ _02910_ _03423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_186_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_246_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09517_ _04543_ _00867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06729_ _02420_ _00202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_168_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_213_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09448_ soc.rom_encoder_0.request_address\[14\] _02520_ _04460_ soc.rom_encoder_0.output_buffer\[11\]
+ _04496_ _04497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XPHY_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_125_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_240_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09379_ soc.spi_video_ram_1.state_sram_clk_counter\[7\] _04445_ _04433_ _04447_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_138_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11410_ _00476_ clknet_leaf_44_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[2\]\[20\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_205_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_181_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11341_ _00407_ clknet_leaf_199_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[27\]\[9\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_193_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11272_ _00338_ clknet_leaf_166_wb_clk_i soc.ram_encoder_0.output_buffer\[18\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_134_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10223_ _05038_ _01078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_152_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_70_wb_clk_i clknet_5_9_0_wb_clk_i clknet_leaf_70_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_10154_ _02485_ _04917_ _04991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_5920 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5931 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5942 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_23_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_66_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5953 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10085_ _04787_ _04938_ _01039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_130_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5964 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_87_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5975 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_212_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5986 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5997 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_236_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_210_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_147_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10987_ _00053_ clknet_leaf_2_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[17\]\[12\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_128_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_128_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_245_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_245_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_230_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_223_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_1242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11608_ _00674_ clknet_leaf_307_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[21\]\[15\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_50_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_191_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11539_ _00605_ clknet_leaf_141_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[25\]\[4\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_128_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_125_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_135_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08750_ soc.spi_video_ram_1.write_fifo.fifo_mem\[24\]\[11\] _02414_ _04087_ _04089_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_85_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05962_ _01852_ _01854_ _01855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XTAP_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_238_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07701_ soc.spi_video_ram_1.write_fifo.fifo_mem\[29\]\[24\] _03347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_6_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08681_ _04031_ _04048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_05893_ _01775_ _01788_ _01789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_65_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_226_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07632_ soc.spi_video_ram_1.current_state\[1\] _02624_ _03279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_4_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07563_ soc.spi_video_ram_1.write_fifo.fifo_mem\[9\]\[13\] _03210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09302_ _04401_ _00793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06514_ _02149_ soc.spi_video_ram_1.write_fifo.fifo_mem\[0\]\[14\] _02290_ _02295_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_07494_ _03139_ soc.spi_video_ram_1.write_fifo.fifo_mem\[14\]\[12\] _03141_ _02646_
+ _03142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_107_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_222_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09233_ _02223_ soc.spi_video_ram_1.write_fifo.fifo_mem\[9\]\[3\] _04360_ _04364_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_167_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06445_ soc.spi_video_ram_1.fifo_in_address\[1\] _02252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xclkbuf_4_15_0_wb_clk_i clknet_3_7_0_wb_clk_i clknet_4_15_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_72_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09164_ soc.video_generator_1.v_count\[2\] _04321_ _04322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06376_ _02206_ _00063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_124_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_120_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08115_ soc.video_generator_1.h_count\[4\] _03717_ _03719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_175_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09095_ _02252_ soc.spi_video_ram_1.write_fifo.fifo_mem\[20\]\[17\] _04270_ _04278_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_11_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_198_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08046_ soc.spi_video_ram_1.write_fifo.fifo_mem\[11\]\[1\] _02393_ _03680_ _03682_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_200_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_131_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_192_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09997_ _04883_ _01007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_103_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_5227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08948_ _04195_ _00645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_4515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_130_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3803 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3814 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_229_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08879_ _04158_ _00613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_91_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_218_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3825 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3836 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_229_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3847 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10910_ soc.spi_video_ram_1.write_fifo.fifo_mem\[8\]\[11\] soc.spi_video_ram_1.fifo_in_data\[11\]
+ _05442_ _05444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_3858 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_211_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3869 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11890_ _00949_ clknet_leaf_25_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[3\]\[16\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10841_ _03354_ _05392_ _05406_ _01328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_71_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_246_1542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_164_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10772_ _03566_ _05358_ _05369_ _01296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_241_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_198_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_212_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_233_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_200_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_1535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_126_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11324_ _00390_ clknet_leaf_231_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[26\]\[21\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_181_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_158_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11255_ _00321_ clknet_leaf_280_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[10\]\[26\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_153_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10206_ _02179_ _04392_ _05029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_84_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_6440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11186_ _00252_ clknet_leaf_58_wb_clk_i soc.spi_video_ram_1.output_buffer\[4\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_6451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_171_1246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_122_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10137_ soc.ram_data_out\[13\] _04928_ _04978_ _04979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5750 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5761 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5772 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_276_wb_clk_i clknet_5_6_0_wb_clk_i clknet_leaf_276_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_94_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5783 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10068_ _04915_ _04923_ _01037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_5794 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_47_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_205_wb_clk_i clknet_5_22_0_wb_clk_i clknet_leaf_205_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_110_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_208_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_63_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_235_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_232_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_204_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_182_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_231_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_188_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06230_ net81 _02112_ net82 vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_15_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_06161_ _01853_ soc.video_generator_1.v_count\[8\] _02054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_176_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_219_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06092_ _01977_ _01981_ _01984_ _01985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_195_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_236_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09920_ soc.rom_encoder_0.initializing_step\[3\] soc.rom_encoder_0.initializing_step\[2\]
+ soc.rom_encoder_0.initializing_step\[1\] _02459_ _04827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_67_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_160_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_193_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09851_ _04752_ _04774_ _00970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_119_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08802_ _04109_ _04117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_86_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09782_ _02262_ soc.spi_video_ram_1.write_fifo.fifo_mem\[3\]\[22\] _04696_ _04721_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_112_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06994_ _02650_ _02653_ _02618_ _02654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_80_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_239_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08733_ soc.spi_video_ram_1.write_fifo.fifo_mem\[24\]\[3\] _02397_ _04076_ _04080_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_05945_ _01837_ _01838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_66_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_227_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08664_ soc.spi_video_ram_1.write_fifo.fifo_mem\[15\]\[5\] _02401_ _04032_ _04038_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_05876_ _01717_ _01772_ _01773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_96_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_241_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07615_ _02582_ _03258_ _03261_ _03262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_1708 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_198_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1719 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_148_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08595_ _02122_ soc.spi_video_ram_1.write_fifo.fifo_mem\[30\]\[1\] _04000_ _04002_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_82_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07546_ soc.spi_video_ram_1.write_fifo.fifo_mem\[18\]\[13\] soc.spi_video_ram_1.write_fifo.fifo_mem\[19\]\[13\]
+ _02651_ _03193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_223_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_201_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07477_ _02901_ _03117_ _03124_ _02970_ _03125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_50_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09216_ _04047_ _04346_ _04354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_52_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06428_ soc.spi_video_ram_1.write_fifo.fifo_mem\[16\]\[11\] _02240_ _02238_ _02241_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_210_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_206_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09147_ _04293_ _04308_ _04309_ _00730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_06359_ _02149_ soc.spi_video_ram_1.write_fifo.fifo_mem\[17\]\[14\] _02193_ _02198_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xclkbuf_5_4_0_wb_clk_i clknet_4_2_0_wb_clk_i clknet_5_4_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_136_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09078_ _02235_ soc.spi_video_ram_1.write_fifo.fifo_mem\[20\]\[9\] _04259_ _04269_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_146_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08029_ _02736_ _03666_ _03667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_122_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_46_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11040_ _00106_ clknet_leaf_205_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[0\]\[7\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_5002 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_89_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5013 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_104_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5024 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5035 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_49_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_5046 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_172_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5057 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_5068 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5079 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_170_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11942_ _01001_ clknet_leaf_159_wb_clk_i soc.ram_encoder_0.input_buffer\[8\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_4378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2910 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2921 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2932 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_217_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2943 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11873_ _00932_ clknet_leaf_165_wb_clk_i net61 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2954 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3699 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2965 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2976 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_214_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2987 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10824_ _02250_ soc.spi_video_ram_1.write_fifo.fifo_mem\[7\]\[16\] _05389_ _05398_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_2998 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_246_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_186_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_213_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10755_ _04050_ _05359_ _05361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_203_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_224_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_199_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_1242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10686_ _02240_ soc.spi_video_ram_1.write_fifo.fifo_mem\[29\]\[11\] _05321_ _05323_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_145_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11307_ _00373_ clknet_leaf_141_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[26\]\[4\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_141_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12287_ _01315_ clknet_leaf_41_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[7\]\[11\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_206_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11238_ _00304_ clknet_leaf_256_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[10\]\[9\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_122_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11169_ _00235_ clknet_leaf_55_wb_clk_i soc.spi_video_ram_1.output_buffer\[21\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_6281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_132_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_95_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_5580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_23_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_110_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05730_ _01628_ _01634_ _01627_ _01635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_212_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_209_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4890 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_223_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05661_ soc.cpu.AReg.data\[11\] soc.cpu.AReg.data\[10\] soc.cpu.AReg.data\[12\] soc.cpu.AReg.data\[5\]
+ _01569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_35_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_149_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07400_ _03021_ soc.spi_video_ram_1.write_fifo.fifo_mem\[11\]\[11\] _02652_ _03049_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_51_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_1702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_75_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08380_ soc.spi_video_ram_1.write_fifo.fifo_mem\[26\]\[18\] _02339_ _03877_ _03886_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_05592_ _01467_ _01501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_205_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07331_ _02696_ soc.spi_video_ram_1.write_fifo.fifo_mem\[9\]\[28\] _02927_ _02981_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_108_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_1749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07262_ _02620_ _02892_ _02912_ _02606_ _02913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_192_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_203_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09001_ _04223_ _00670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_118_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06213_ _01469_ soc.spi_video_ram_1.output_buffer\[1\] _01492_ _02099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_30_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_192_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07193_ _01419_ _02846_ _02847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_118_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06144_ _01849_ _01939_ _01940_ _02037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_133_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_191_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06075_ soc.video_generator_1.h_count\[1\] soc.display_clks_before_active\[0\] _01968_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_117_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09903_ _04809_ _04813_ _04814_ _04254_ _00982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_63_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_198_wb_clk_i clknet_5_25_0_wb_clk_i clknet_leaf_198_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_67_1282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_154_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_63_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_236_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09834_ _04742_ _04761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
Xclkbuf_leaf_127_wb_clk_i clknet_5_13_0_wb_clk_i clknet_leaf_127_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_63_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_58_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_150_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09765_ _04712_ _00946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06977_ soc.spi_video_ram_1.write_fifo.fifo_mem\[8\]\[1\] soc.spi_video_ram_1.write_fifo.fifo_mem\[9\]\[1\]
+ soc.spi_video_ram_1.write_fifo.fifo_mem\[10\]\[1\] soc.spi_video_ram_1.write_fifo.fifo_mem\[11\]\[1\]
+ _02635_ _02636_ _02637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_246_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_189_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_230_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08716_ _04069_ _04048_ _04070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_210_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05928_ _01702_ _01821_ _01822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_55_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09696_ _04639_ soc.rom_loader.current_address\[10\] _04665_ _04666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_27_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_148_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08647_ _04028_ _00511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_55_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_199_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05859_ _01670_ soc.cpu.ALU.x\[10\] _01757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_81_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_08578_ _02167_ soc.spi_video_ram_1.write_fifo.fifo_mem\[2\]\[23\] _03966_ _03992_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_39_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_242_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_186_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_126_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07529_ _02700_ soc.spi_video_ram_1.write_fifo.fifo_mem\[6\]\[26\] _03176_ _02577_
+ _03177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_70_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10540_ soc.ram_encoder_0.address\[11\] soc.cpu.AReg.data\[11\] _05227_ _05240_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_10_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_211_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_168_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_241_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_196_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10471_ soc.cpu.PC.in\[6\] _05188_ _05173_ _05192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_6_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12210_ _01238_ clknet_leaf_241_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[19\]\[21\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_157_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12141_ _01169_ net88 soc.cpu.PC.REG.data\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_123_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_155_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12072_ _01115_ clknet_leaf_109_wb_clk_i soc.rom_loader.current_address\[12\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_89_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_172_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11023_ _00089_ clknet_leaf_67_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[16\]\[19\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_81_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4120 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4131 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_77_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4142 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4153 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4164 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4175 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_4186 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_205_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11925_ _00984_ clknet_leaf_86_wb_clk_i soc.rom_encoder_0.initializing_step\[0\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2740 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2751 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_221_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2762 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2773 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11856_ _00915_ clknet_leaf_107_wb_clk_i soc.rom_encoder_0.request_address\[1\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_33_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2784 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2795 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_207_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10807_ _02235_ soc.spi_video_ram_1.write_fifo.fifo_mem\[7\]\[9\] _05378_ _05388_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_57_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_60_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11787_ _00848_ clknet_leaf_102_wb_clk_i soc.rom_encoder_0.output_buffer\[18\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_13_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10738_ soc.spi_video_ram_1.write_fifo.fifo_mem\[31\]\[6\] soc.spi_video_ram_1.fifo_in_data\[6\]
+ _05344_ _05351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_119_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_9_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_242_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_31_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10669_ _02223_ soc.spi_video_ram_1.write_fifo.fifo_mem\[29\]\[3\] _05310_ _05314_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_51_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_86_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_220_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12339_ _01367_ clknet_leaf_26_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[8\]\[18\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_47_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_233_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_291_wb_clk_i clknet_5_5_0_wb_clk_i clknet_leaf_291_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_64_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_214_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_155_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06900_ _02555_ _02563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_151_1403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_leaf_220_wb_clk_i clknet_5_21_0_wb_clk_i clknet_leaf_220_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_64_1477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07880_ _01885_ _02625_ _03523_ _03524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06831_ _02505_ _02506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_3_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_231_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09550_ _04243_ _04252_ _04253_ _00880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_06762_ soc.rom_encoder_0.output_bits_left\[4\] _02440_ _02441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_149_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08501_ _03951_ _00442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05713_ soc.cpu.AReg.data\[2\] _01619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_236_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09481_ _01485_ _04521_ _04523_ _04519_ _00851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_64_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06693_ soc.spi_video_ram_1.write_fifo.fifo_mem\[14\]\[3\] _02397_ _02391_ _02398_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_91_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08432_ soc.spi_video_ram_1.write_fifo.fifo_mem\[27\]\[13\] _02244_ _03910_ _03914_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_197_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05644_ soc.cpu.instruction\[15\] _01552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_52_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_224_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_184_1278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_211_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_168_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_162_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08363_ _03864_ _03877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_05575_ _01468_ soc.spi_video_ram_1.output_buffer\[6\] _01477_ soc.spi_video_ram_1.output_buffer\[7\]
+ _01484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_108_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07314_ _02573_ soc.spi_video_ram_1.write_fifo.fifo_mem\[29\]\[10\] _02964_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_165_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08294_ _03839_ _00347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_109_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07245_ soc.spi_video_ram_1.write_fifo.fifo_mem\[28\]\[9\] soc.spi_video_ram_1.write_fifo.fifo_mem\[29\]\[9\]
+ soc.spi_video_ram_1.write_fifo.fifo_mem\[30\]\[9\] soc.spi_video_ram_1.write_fifo.fifo_mem\[31\]\[9\]
+ _02893_ _02895_ _02896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_197_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_191_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_180_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07176_ soc.spi_video_ram_1.write_fifo.fifo_mem\[28\]\[6\] soc.spi_video_ram_1.write_fifo.fifo_mem\[29\]\[6\]
+ soc.spi_video_ram_1.write_fifo.fifo_mem\[30\]\[6\] soc.spi_video_ram_1.write_fifo.fifo_mem\[31\]\[6\]
+ _02680_ _02722_ _02830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_173_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06127_ _02016_ _02019_ _01986_ _02020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_30_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_308_wb_clk_i clknet_5_1_0_wb_clk_i clknet_leaf_308_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_105_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06058_ _01949_ _01844_ _01947_ _01951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_133_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_1544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_87_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_87_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09817_ _01396_ _04747_ _00963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_234_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09748_ _04703_ _00938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_228_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2003 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2014 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2025 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_210_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09679_ _04653_ _00919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_54_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2036 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2047 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_203_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_95_wb_clk_i clknet_5_11_0_wb_clk_i clknet_leaf_95_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_11710_ _00771_ clknet_leaf_2_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[9\]\[12\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2058 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2069 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_226_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_24_wb_clk_i clknet_5_8_0_wb_clk_i clknet_leaf_24_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_11641_ _00702_ clknet_leaf_256_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[20\]\[9\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_35_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_146_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_204_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_168_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11572_ _00638_ clknet_leaf_208_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[22\]\[8\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_122_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput19 la_data_in[10] net19 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_10523_ _01619_ _05228_ _05231_ _01185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_183_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_171_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xcaravel_hack_soc_210 wbs_dat_o[18] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_10454_ soc.cpu.PC.in\[2\] _05172_ _05173_ _05179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_87_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xcaravel_hack_soc_221 wbs_dat_o[29] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_237_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10385_ _02235_ soc.spi_video_ram_1.write_fifo.fifo_mem\[6\]\[9\] _05124_ _05134_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_100_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12124_ _01152_ clknet_leaf_75_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[6\]\[16\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_215_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_238_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12055_ net33 clknet_opt_2_0_wb_clk_i soc.rom_encoder_0.data_out\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_152_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11006_ _00072_ clknet_leaf_197_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[16\]\[2\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_24_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_218_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_59_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11908_ _00967_ clknet_leaf_127_wb_clk_i soc.cpu.instruction\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_34_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_206_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11839_ _00898_ clknet_leaf_102_wb_clk_i soc.rom_encoder_0.request_data_out\[0\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_21_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1891 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07030_ _02688_ _02689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_173_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_162_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_61_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_200_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_192_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_244_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08981_ soc.spi_video_ram_1.write_fifo.fifo_mem\[21\]\[2\] _02395_ _04210_ _04213_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_244_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07932_ _03574_ _00250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_138_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_228_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07863_ _02952_ _03503_ _03506_ _03507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_69_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_244_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_151_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06814_ _02481_ _02482_ _02490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09602_ soc.rom_encoder_0.input_buffer\[8\] _04603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_99_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_216_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07794_ soc.spi_video_ram_1.write_fifo.fifo_mem\[24\]\[23\] soc.spi_video_ram_1.write_fifo.fifo_mem\[25\]\[23\]
+ soc.spi_video_ram_1.write_fifo.fifo_mem\[26\]\[23\] soc.spi_video_ram_1.write_fifo.fifo_mem\[27\]\[23\]
+ _02903_ _02904_ _03439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_09533_ _01444_ _04552_ _04554_ _00872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_243_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06745_ _02428_ _00210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_36_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_129_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_240_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09464_ _02443_ _04509_ _04510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06676_ _02175_ soc.spi_video_ram_1.write_fifo.fifo_mem\[12\]\[27\] _02356_ _02386_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_227_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_149_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_169_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_149_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08415_ soc.spi_video_ram_1.write_fifo.fifo_mem\[27\]\[5\] _02401_ _03899_ _03905_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_184_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05627_ _01501_ _01534_ _01535_ _01536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_09395_ _02061_ _04454_ _04456_ _00832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_196_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_205_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08346_ _03868_ _00370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_149_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05558_ _01461_ _01467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_127_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_165_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08277_ _03829_ _03830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_165_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05489_ soc.spi_video_ram_1.write_fifo.read_pointer\[3\] _01403_ _01404_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_123_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07228_ _02606_ _02879_ _02880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_leaf_142_wb_clk_i clknet_5_25_0_wb_clk_i clknet_leaf_142_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_07159_ _02583_ _02813_ _02640_ _02814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_69_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_161_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_234_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10170_ soc.ram_encoder_0.toggled_sram_sck _02492_ _05003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_154_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_235_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_41_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_245_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_16_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_245_1448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_182_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_230_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_167_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11624_ _00690_ clknet_leaf_32_wb_clk_i _00002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_169_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_184_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11555_ _00621_ clknet_leaf_263_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[25\]\[20\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_32_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_11_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_102_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_10_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10506_ net90 _05218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_155_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11486_ _00552_ clknet_leaf_201_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[24\]\[9\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_13_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10437_ _01779_ _01819_ _05163_ _05164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_100_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_151_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10368_ _05125_ _01136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_83_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12107_ _01135_ net85 soc.cpu.ALU.x\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_239_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10299_ soc.rom_loader.current_address\[6\] _05082_ _05083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_214_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_12038_ _01097_ clknet_leaf_295_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[5\]\[26\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_78_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_226_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_211_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_225_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_81_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06530_ _02165_ soc.spi_video_ram_1.write_fifo.fifo_mem\[0\]\[22\] _02278_ _02303_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_222_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_185_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3090 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_209_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06461_ soc.spi_video_ram_1.write_fifo.fifo_mem\[16\]\[22\] _02262_ _02216_ _02263_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_221_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08200_ _02460_ _03764_ _03769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_33_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09180_ _02034_ _04325_ _04333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06392_ _02215_ _02216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_30_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08131_ _02116_ _03677_ _03729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_120_1508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_198_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_200_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08062_ soc.spi_video_ram_1.write_fifo.fifo_mem\[11\]\[9\] _02409_ _03680_ _03690_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_179_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07013_ _02624_ _02671_ _02672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_190_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_235_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_5409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_130_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08964_ _04203_ _00653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_102_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_229_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4708 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07915_ _02613_ _03557_ _03558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_124_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4719 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08895_ _04166_ _00621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_130_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_245_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07846_ soc.spi_video_ram_1.write_fifo.fifo_mem\[24\]\[22\] soc.spi_video_ram_1.write_fifo.fifo_mem\[25\]\[22\]
+ soc.spi_video_ram_1.write_fifo.fifo_mem\[26\]\[22\] soc.spi_video_ram_1.write_fifo.fifo_mem\[27\]\[22\]
+ _02893_ _02895_ _03490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_217_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07777_ _02588_ _03418_ _03421_ _03422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_99_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_37_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_56_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09516_ _02270_ soc.cpu.AReg.data\[10\] _01459_ _04543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06728_ soc.spi_video_ram_1.write_fifo.fifo_mem\[14\]\[16\] _02335_ _02412_ _02420_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_25_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_246_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_212_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09447_ soc.rom_encoder_0.request_data_out\[7\] _03767_ _04496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XPHY_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_242_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_164_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06659_ _02377_ _00175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_197_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_240_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_200_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09378_ _04445_ _04446_ _00824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_138_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_162_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08329_ _03857_ _00364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_71_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_166_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11340_ _00406_ clknet_leaf_184_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[27\]\[8\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_126_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_192_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_166_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_197_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11271_ _00337_ clknet_leaf_166_wb_clk_i soc.ram_encoder_0.output_buffer\[17\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_106_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_238_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10222_ _02231_ soc.spi_video_ram_1.write_fifo.fifo_mem\[5\]\[7\] _05030_ _05038_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_88_1594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10153_ _04990_ _01055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_5910 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_5921 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_47_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5932 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5943 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10084_ soc.ram_data_out\[1\] _04927_ _04937_ _04938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_5954 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5965 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5976 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_208_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5987 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5998 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_207_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_204_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_16_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10986_ _00052_ clknet_leaf_37_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[17\]\[11\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_128_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_231_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_188_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_203_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_15_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11607_ _00673_ clknet_leaf_308_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[21\]\[14\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_157_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11538_ _00604_ clknet_leaf_142_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[25\]\[3\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_144_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_183_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11469_ _00535_ clknet_leaf_283_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[15\]\[21\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_48_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_215_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05961_ soc.video_generator_1.v_count\[3\] _01851_ _01850_ _01853_ _01854_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_24_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_230_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07700_ _02590_ soc.spi_video_ram_1.write_fifo.fifo_mem\[30\]\[24\] _03345_ _02576_
+ _03346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_227_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_152_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_152_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08680_ soc.spi_video_ram_1.fifo_in_data\[12\] _04047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_05892_ _01762_ _01776_ _01788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_96_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07631_ _02918_ _03254_ _03277_ _03278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_66_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07562_ _02922_ soc.spi_video_ram_1.write_fifo.fifo_mem\[11\]\[13\] _02647_ _03209_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_94_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_228_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09301_ _02227_ soc.spi_video_ram_1.write_fifo.fifo_mem\[4\]\[5\] _04395_ _04401_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06513_ _02294_ _00112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07493_ _02644_ _03140_ _03141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_34_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09232_ _04363_ _00761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06444_ _02251_ _00086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_206_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_181_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_241_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_222_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_163_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09163_ _04317_ _04320_ _04321_ _00734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_06375_ _02165_ soc.spi_video_ram_1.write_fifo.fifo_mem\[17\]\[22\] _02181_ _02206_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_08114_ _03713_ _03717_ _03718_ _00288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_119_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09094_ _04277_ _00709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_135_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_190_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08045_ _03681_ _00256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_163_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_239_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09996_ soc.ram_encoder_0.request_data_out\[1\] soc.ram_encoder_0.data_out\[1\] _04880_
+ _04883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_89_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_170_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08947_ soc.spi_video_ram_1.write_fifo.fifo_mem\[22\]\[15\] _04054_ _04189_ _04195_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_4516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3804 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3815 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08878_ soc.spi_video_ram_1.write_fifo.fifo_mem\[25\]\[12\] _04047_ _04155_ _04158_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_3826 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3837 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_244_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07829_ soc.video_generator_1.v_count\[2\] _01897_ _03474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_3848 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3859 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10840_ soc.spi_video_ram_1.fifo_in_address\[8\] _05393_ _05406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_213_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10771_ _04061_ _05359_ _05369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_92_1749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_240_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_13_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_201_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_226_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_205_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_220_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_193_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_165_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11323_ _00389_ clknet_leaf_52_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[26\]\[20\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_154_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_107_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11254_ _00320_ clknet_leaf_236_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[10\]\[25\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_141_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_45_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10205_ _05017_ _05028_ _01070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_136_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_218_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11185_ _00251_ clknet_leaf_59_wb_clk_i soc.spi_video_ram_1.output_buffer\[5\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_45_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_68_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10136_ _04867_ _04947_ _04948_ _04977_ _04978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_6474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_122_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5740 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5751 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5762 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_212_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_209_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5773 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10067_ _04918_ _01059_ _04923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_5784 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5795 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_236_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_149_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_62_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_245_wb_clk_i clknet_5_17_0_wb_clk_i clknet_leaf_245_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_189_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10969_ _00035_ clknet_leaf_234_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[18\]\[23\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_223_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06160_ soc.hack_wait_clocks\[1\] soc.hack_wait_clocks\[0\] _01452_ _01453_ _02053_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_141_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06091_ _01976_ _01983_ _01984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_144_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_236_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_158_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09850_ _01669_ _04740_ _04773_ _04774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08801_ _04116_ _00577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_98_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09781_ _04720_ _00954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06993_ soc.spi_video_ram_1.write_fifo.fifo_mem\[4\]\[1\] soc.spi_video_ram_1.write_fifo.fifo_mem\[5\]\[1\]
+ soc.spi_video_ram_1.write_fifo.fifo_mem\[6\]\[1\] soc.spi_video_ram_1.write_fifo.fifo_mem\[7\]\[1\]
+ _02651_ _02652_ _02653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_85_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05944_ soc.video_generator_1.h_count\[5\] soc.video_generator_1.h_count\[6\] soc.video_generator_1.h_count\[7\]
+ _01837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_6_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08732_ _04079_ _00545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_61_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_187_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08663_ _04037_ _00518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_226_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05875_ _01618_ soc.cpu.AReg.data\[11\] _01718_ soc.ram_data_out\[11\] _01772_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_187_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_148_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07614_ _02971_ soc.spi_video_ram_1.write_fifo.fifo_mem\[6\]\[25\] _03260_ _02838_
+ _03261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_1709 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08594_ _04001_ _00485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_242_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_1413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07545_ _03041_ _03188_ _03191_ _02570_ _03192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_243_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_241_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_222_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07476_ _02642_ _03120_ _03123_ _03124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_09215_ _04341_ _01779_ _04353_ _00754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06427_ soc.spi_video_ram_1.fifo_in_data\[11\] _02240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_72_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_72_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09146_ soc.spi_video_ram_1.state_counter\[8\] _04306_ _04309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06358_ _02197_ _00054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_202_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_194_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_33_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_147_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_198_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09077_ _04268_ _00701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_205_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06289_ _02154_ _00028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_120_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_120_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_200_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08028_ soc.spi_video_ram_1.write_fifo.fifo_mem\[24\]\[16\] soc.spi_video_ram_1.write_fifo.fifo_mem\[25\]\[16\]
+ soc.spi_video_ram_1.write_fifo.fifo_mem\[26\]\[16\] soc.spi_video_ram_1.write_fifo.fifo_mem\[27\]\[16\]
+ _02701_ _02737_ _03666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
Xclkbuf_leaf_49_wb_clk_i clknet_5_13_0_wb_clk_i clknet_leaf_49_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_155_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_81_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_5003 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_235_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5014 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5025 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5036 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09979_ soc.ram_encoder_0.input_buffer\[6\] _04847_ _04248_ _04870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_162_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5047 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_118_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5058 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5069 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_213_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_218_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11941_ _01000_ clknet_leaf_159_wb_clk_i soc.ram_encoder_0.input_buffer\[7\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_4379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_176_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_44_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2900 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2911 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2922 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2933 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11872_ _00931_ clknet_leaf_165_wb_clk_i net60 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2944 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2955 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2966 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2977 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10823_ _03416_ _05392_ _05397_ _01319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_60_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2988 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2999 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_241_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_198_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_242_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10754_ _03121_ _05358_ _05360_ _01287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_57_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10685_ _05322_ _01256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_200_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11306_ _00372_ clknet_leaf_142_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[26\]\[3\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_154_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12286_ _01314_ clknet_leaf_13_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[7\]\[10\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_153_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11237_ _00303_ clknet_leaf_190_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[10\]\[8\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_155_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_190_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11168_ _00234_ clknet_leaf_56_wb_clk_i soc.spi_video_ram_1.output_buffer\[22\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_110_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10119_ soc.ram_encoder_0.request_data_out\[9\] _04929_ _04965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_110_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11099_ _00165_ clknet_leaf_175_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[12\]\[8\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_5581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_222_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_208_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4880 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4891 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05660_ soc.cpu.AReg.data\[4\] soc.cpu.AReg.data\[7\] soc.cpu.AReg.data\[6\] _01568_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_63_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_224_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_188_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05591_ _01460_ _01462_ _01466_ _01499_ _01500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_223_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_204_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07330_ _02744_ soc.spi_video_ram_1.write_fifo.fifo_mem\[8\]\[28\] _02980_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_177_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_182_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_220_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_188_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07261_ _02897_ _02899_ _02906_ _02911_ _02567_ _02912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_73_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09000_ soc.spi_video_ram_1.write_fifo.fifo_mem\[21\]\[11\] _02414_ _04221_ _04223_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_118_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06212_ _02097_ _02098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_121_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_176_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07192_ _02623_ _02624_ _02846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_157_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_185_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06143_ soc.video_generator_1.v_count\[1\] _01856_ _01897_ _02035_ _02036_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_219_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_201_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06074_ _01945_ _01963_ _01966_ _01967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
X_09902_ _02435_ _04809_ _04814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_193_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09833_ _04752_ _04760_ _00966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_141_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09764_ _02244_ soc.spi_video_ram_1.write_fifo.fifo_mem\[3\]\[13\] _04708_ _04712_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06976_ _02592_ _02636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_246_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_167_wb_clk_i clknet_5_30_0_wb_clk_i clknet_leaf_167_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_132_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08715_ soc.spi_video_ram_1.fifo_in_address\[9\] _04069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_05927_ _01670_ soc.cpu.ALU.x\[14\] _01821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_100_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_227_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09695_ _04639_ _04664_ _04665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_26_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05858_ _01745_ _01755_ _01756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_27_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08646_ _02173_ soc.spi_video_ram_1.write_fifo.fifo_mem\[30\]\[26\] _03999_ _04028_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XPHY_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_35 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05789_ _01663_ _01690_ _01691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XPHY_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_08577_ _03991_ _00478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_35_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_223_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07528_ _02574_ _03175_ _03176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_243_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07459_ _01940_ _03106_ _03107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_168_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_210_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10470_ soc.cpu.PC.REG.data\[6\] _05190_ _05191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_52_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09129_ _04294_ _04296_ _04297_ _00724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_100_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12140_ _01168_ net88 soc.cpu.PC.REG.data\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_139_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_191_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_151_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_190_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_12071_ _01114_ clknet_leaf_110_wb_clk_i soc.rom_loader.current_address\[11\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_194_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_151_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11022_ _00088_ clknet_leaf_75_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[16\]\[18\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_172_1353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_172_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4110 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4121 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4132 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4143 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4154 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4165 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_185_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4176 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_3431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4187 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11924_ _00983_ clknet_leaf_98_wb_clk_i soc.rom_encoder_0.current_state\[2\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XTAP_3464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_206_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_166_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2730 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2741 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_209_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2752 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2763 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11855_ _00914_ clknet_leaf_92_wb_clk_i soc.rom_encoder_0.request_address\[0\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_60_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2774 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2785 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_205_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2796 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10806_ _05387_ _01312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_246_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_199_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11786_ _00847_ clknet_leaf_104_wb_clk_i soc.rom_encoder_0.output_buffer\[17\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_202_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_183_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10737_ _05350_ _01280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_186_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_201_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10668_ _05313_ _01248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_127_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10599_ _01445_ _02117_ _05276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_182_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12338_ _01366_ clknet_leaf_24_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[8\]\[17\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_177_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_5_30_0_wb_clk_i clknet_4_15_0_wb_clk_i clknet_5_30_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_12269_ _01297_ clknet_leaf_268_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[31\]\[22\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_68_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_233_1726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06830_ _02484_ _02503_ _02504_ _02505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XTAP_6090 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_95_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06761_ _02439_ soc.rom_encoder_0.output_bits_left\[2\] _02440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_37_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_260_wb_clk_i clknet_5_18_0_wb_clk_i clknet_leaf_260_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_114_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_209_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05712_ _01563_ _01618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_08500_ _02151_ soc.spi_video_ram_1.write_fifo.fifo_mem\[28\]\[15\] _03945_ _03951_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_64_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06692_ soc.spi_video_ram_1.fifo_in_data\[3\] _02397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_09480_ _01501_ _04521_ _01469_ _04523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_149_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_149_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05643_ _01551_ net70 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_08431_ _03913_ _00410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_64_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_205_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08362_ _03876_ _00378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_177_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05574_ _01467_ soc.spi_video_ram_1.output_buffer\[4\] _01477_ soc.spi_video_ram_1.output_buffer\[5\]
+ _01483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_177_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_32_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_189_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07313_ _02763_ soc.spi_video_ram_1.write_fifo.fifo_mem\[30\]\[10\] _02592_ _02963_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_71_1438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08293_ _02134_ soc.spi_video_ram_1.write_fifo.fifo_mem\[1\]\[7\] _03831_ _03839_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_192_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07244_ _02894_ _02895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_30_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07175_ _02767_ _02828_ _02829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_145_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06126_ _01987_ _02017_ _02018_ _01989_ _02019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_156_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_191_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_172_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06057_ _01844_ _01947_ _01949_ _01950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_47_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_207_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_236_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_154_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09816_ soc.cpu.DMuxJMP.sel\[0\] _04740_ _04746_ _04747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_47_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_214_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09747_ _02227_ soc.spi_video_ram_1.write_fifo.fifo_mem\[3\]\[5\] _04697_ _04703_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06959_ _00004_ _02620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_27_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2004 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2015 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_167_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09678_ _04652_ soc.rom_encoder_0.request_address\[5\] _04632_ _04653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_2026 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_199_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2037 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2048 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2059 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08629_ _04019_ _00502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_188_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_242_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11640_ _00701_ clknet_leaf_208_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[20\]\[8\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_74_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_11_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11571_ _00637_ clknet_leaf_194_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[22\]\[7\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_156_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_211_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_168_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_64_wb_clk_i clknet_5_12_0_wb_clk_i clknet_leaf_64_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_10522_ soc.ram_encoder_0.address\[2\] _05228_ _05231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_182_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xcaravel_hack_soc_200 wbs_dat_o[8] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_10453_ soc.cpu.PC.REG.data\[2\] _05177_ _05178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_100_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xcaravel_hack_soc_211 wbs_dat_o[19] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_164_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xcaravel_hack_soc_222 wbs_dat_o[30] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_202_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10384_ _05133_ _01144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_123_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_174_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_139_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12123_ _01151_ clknet_leaf_316_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[6\]\[15\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_2_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12054_ net32 clknet_leaf_108_wb_clk_i soc.rom_encoder_0.data_out\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_85_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_133_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11005_ _00071_ clknet_leaf_218_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[16\]\[1\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_42_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_238_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11907_ _00966_ clknet_leaf_121_wb_clk_i soc.cpu.instruction\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_234_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_146_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_181_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11838_ _00897_ clknet_leaf_101_wb_clk_i soc.rom_encoder_0.request_write vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_159_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1870 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1881 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1892 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_226_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11769_ _00830_ clknet_leaf_60_wb_clk_i net68 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_174_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_187_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_174_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_1471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_220_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_177_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_154_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08980_ _04212_ _00660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_69_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_29_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07931_ soc.spi_video_ram_1.output_buffer\[6\] _02882_ _03573_ _03574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_68_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07862_ _03047_ soc.spi_video_ram_1.write_fifo.fifo_mem\[4\]\[22\] _03505_ _03024_
+ _03506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_99_1316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09601_ _04600_ _04585_ _04602_ _00892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_111_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06813_ _02479_ _02488_ _02489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_231_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07793_ _02618_ _03437_ _03438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_228_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09532_ _01444_ _04552_ _04553_ _04554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_37_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06744_ soc.spi_video_ram_1.write_fifo.fifo_mem\[14\]\[24\] _02266_ _02390_ _02428_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_25_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_97_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09463_ soc.rom_encoder_0.output_buffer\[14\] _02463_ _02464_ soc.rom_encoder_0.request_data_out\[10\]
+ _04509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_06675_ _02385_ _00183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_197_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_224_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_08414_ _03904_ _00402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05626_ _01467_ soc.spi_video_ram_1.output_buffer\[21\] _01535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09394_ net10 _04454_ _04456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_184_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_244_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_240_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08345_ soc.spi_video_ram_1.write_fifo.fifo_mem\[26\]\[1\] _02393_ _03866_ _03868_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_05557_ _01462_ _01465_ _01466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_71_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_193_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08276_ _02179_ _02276_ _03829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_164_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05488_ soc.spi_video_ram_1.write_fifo.write_pointer\[3\] _01403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_197_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07227_ _02872_ _02874_ _02876_ _02878_ _02620_ _02879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_180_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_153_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07158_ soc.spi_video_ram_1.write_fifo.fifo_mem\[24\]\[5\] soc.spi_video_ram_1.write_fifo.fifo_mem\[25\]\[5\]
+ soc.spi_video_ram_1.write_fifo.fifo_mem\[26\]\[5\] soc.spi_video_ram_1.write_fifo.fifo_mem\[27\]\[5\]
+ _02635_ _02636_ _02813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_49_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_105_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06109_ _01922_ _01979_ _01985_ _02001_ _02002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_161_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07089_ _02697_ soc.spi_video_ram_1.write_fifo.fifo_mem\[7\]\[3\] _02745_ _02723_
+ _02746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_65_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_1353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_111_wb_clk_i clknet_opt_3_0_wb_clk_i clknet_leaf_111_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_134_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_232_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_234_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_21_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_210_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_95_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_216_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_1438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_187_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_223_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_204_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_169_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_145_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11623_ _00689_ clknet_leaf_47_wb_clk_i _00001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_169_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_223_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_156_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11554_ _00620_ clknet_leaf_35_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[25\]\[19\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_183_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10505_ _05172_ _05216_ _05217_ _01180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_239_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11485_ _00551_ clknet_leaf_180_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[24\]\[8\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_221_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_171_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10436_ _05157_ _05158_ _05159_ _05162_ _05163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_139_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_171_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10367_ _02213_ soc.spi_video_ram_1.write_fifo.fifo_mem\[6\]\[0\] _05124_ _05125_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_174_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_170_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12106_ _01134_ net85 soc.cpu.ALU.x\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10298_ _05071_ _05081_ _05082_ _01108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XTAP_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_152_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12037_ _01096_ clknet_leaf_289_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[5\]\[25\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_66_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_239_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_187_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_230_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_240_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3080 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_179_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3091 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_206_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06460_ soc.spi_video_ram_1.fifo_in_address\[6\] _02262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_59_1388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_146_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_107_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_222_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06391_ _02117_ _02214_ _02215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_175_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08130_ _03713_ _03728_ _00294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_175_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08061_ _03689_ _00264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_70_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_88_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07012_ _02630_ _02631_ _02671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_162_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_239_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_192_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_200_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_216_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08963_ soc.spi_video_ram_1.write_fifo.fifo_mem\[22\]\[23\] _04065_ _04177_ _04203_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_29_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07914_ soc.spi_video_ram_1.write_fifo.fifo_mem\[21\]\[21\] _03557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_116_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4709 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08894_ soc.spi_video_ram_1.write_fifo.fifo_mem\[25\]\[20\] _02343_ _04143_ _04166_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_84_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07845_ _02602_ _03488_ _03489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_96_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_216_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_57_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_229_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07776_ _02924_ soc.spi_video_ram_1.write_fifo.fifo_mem\[4\]\[15\] _03420_ _02927_
+ _03421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_77_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_1714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09515_ _04542_ _00866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06727_ _02419_ _00201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_227_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09446_ _04473_ _04494_ _04495_ _00844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_169_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06658_ _02157_ soc.spi_video_ram_1.write_fifo.fifo_mem\[12\]\[18\] _02368_ _02377_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XPHY_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_205_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05609_ _01470_ _01518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09377_ soc.spi_video_ram_1.state_sram_clk_counter\[6\] _04443_ _04433_ _04446_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_36_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06589_ soc.spi_video_ram_1.write_fifo.fifo_mem\[13\]\[17\] _02337_ _02328_ _02338_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_142_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08328_ _02169_ soc.spi_video_ram_1.write_fifo.fifo_mem\[1\]\[24\] _03830_ _03857_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_32_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_165_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_20_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_240_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08259_ soc.ram_encoder_0.request_write _03816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_166_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_20_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_181_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_153_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11270_ _00336_ clknet_leaf_167_wb_clk_i soc.ram_encoder_0.output_buffer\[16\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_118_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10221_ _05037_ _01077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_49_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10152_ soc.ram_encoder_0.sram_sio_oe _04878_ _04880_ _01395_ _04990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_161_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_239_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5900 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_5911 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5922 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5933 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10083_ _04928_ _04935_ _04936_ _04937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_5944 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5955 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_130_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5966 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_181_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5977 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5988 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5999 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_235_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_74_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_245_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_222_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10985_ _00051_ clknet_leaf_13_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[17\]\[10\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_182_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_204_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_176_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11606_ _00672_ clknet_leaf_41_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[21\]\[13\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_128_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11537_ _00603_ clknet_leaf_196_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[25\]\[2\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_144_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11468_ _00534_ clknet_leaf_50_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[15\]\[20\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_143_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_193_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10419_ _05151_ _01161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_125_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11399_ _00465_ clknet_leaf_249_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[2\]\[9\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_217_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05960_ soc.video_generator_1.v_count\[9\] _01853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XTAP_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05891_ _01729_ _01746_ _01787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_17_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07630_ _02656_ _03263_ _03276_ _03277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_54_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_93_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07561_ _02920_ soc.spi_video_ram_1.write_fifo.fifo_mem\[10\]\[13\] _03208_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_241_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_185_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09300_ _04400_ _00792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06512_ _02147_ soc.spi_video_ram_1.write_fifo.fifo_mem\[0\]\[13\] _02290_ _02294_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_94_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_224_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07492_ soc.spi_video_ram_1.write_fifo.fifo_mem\[15\]\[12\] _03140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_80_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_221_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_210_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09231_ _02221_ soc.spi_video_ram_1.write_fifo.fifo_mem\[9\]\[2\] _04360_ _04363_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_181_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_22_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06443_ soc.spi_video_ram_1.write_fifo.fifo_mem\[16\]\[16\] _02250_ _02238_ _02251_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_72_1352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_194_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09162_ soc.video_generator_1.v_count\[1\] _04313_ _04321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_9_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06374_ _02205_ _00062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_147_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_198_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_241_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08113_ soc.video_generator_1.h_count\[2\] _03715_ soc.video_generator_1.h_count\[3\]
+ _03718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_163_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09093_ _02250_ soc.spi_video_ram_1.write_fifo.fifo_mem\[20\]\[16\] _04270_ _04277_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_163_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08044_ soc.spi_video_ram_1.write_fifo.fifo_mem\[11\]\[0\] _02310_ _03680_ _03681_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_235_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_172_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09995_ _04882_ _01006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_130_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08946_ _04194_ _00644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_103_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_4528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_245_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_3805 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08877_ _04157_ _00612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_111_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_217_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3816 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3827 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3838 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07828_ _03425_ _03472_ _03279_ _03473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_84_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3849 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_233_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_204_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07759_ soc.spi_video_ram_1.write_fifo.fifo_mem\[15\]\[15\] _03404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_72_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_198_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_129_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10770_ _05368_ _01295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_246_1577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_164_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_197_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09429_ soc.rom_encoder_0.output_buffer\[10\] _04479_ _04483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_200_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_201_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_219_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_1559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11322_ _00388_ clknet_leaf_35_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[26\]\[19\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_197_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_158_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_10_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_88_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11253_ _00319_ clknet_leaf_304_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[10\]\[24\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_4_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10204_ soc.hack_clock_0.counter\[6\] _05027_ _05028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_6420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11184_ _00250_ clknet_leaf_56_wb_clk_i soc.spi_video_ram_1.output_buffer\[6\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_6431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_122_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10135_ soc.ram_encoder_0.request_data_out\[13\] _04929_ _04977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_136_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5730 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5741 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_125_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5752 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5763 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10066_ soc.ram_encoder_0.initializing_step\[0\] _04919_ _04922_ _01378_ _01059_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XTAP_5774 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_134_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_5785 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5796 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_223_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_189_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_188_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10968_ _00034_ clknet_leaf_252_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[18\]\[22\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_62_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_225_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_203_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10899_ soc.spi_video_ram_1.write_fifo.fifo_mem\[8\]\[6\] soc.spi_video_ram_1.fifo_in_data\[6\]
+ _05431_ _05438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_176_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_285_wb_clk_i clknet_5_5_0_wb_clk_i clknet_leaf_285_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_129_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_141_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_214_wb_clk_i clknet_5_20_0_wb_clk_i clknet_leaf_214_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_145_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06090_ _01967_ _01982_ _01983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_195_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_172_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_236_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_154_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08800_ _02130_ soc.spi_video_ram_1.write_fifo.fifo_mem\[23\]\[5\] _04110_ _04116_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09780_ _02260_ soc.spi_video_ram_1.write_fifo.fifo_mem\[3\]\[21\] _04696_ _04720_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06992_ _02592_ _02652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_246_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_230_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08731_ soc.spi_video_ram_1.write_fifo.fifo_mem\[24\]\[2\] _02395_ _04076_ _04079_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_227_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_152_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05943_ soc.video_generator_1.h_count\[5\] _01836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_26_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08662_ soc.spi_video_ram_1.write_fifo.fifo_mem\[15\]\[4\] _02399_ _04032_ _04037_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_187_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_05874_ _01702_ _01770_ _01771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_215_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07613_ _02763_ _03259_ _03260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_81_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_187_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_54_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08593_ _02113_ soc.spi_video_ram_1.write_fifo.fifo_mem\[30\]\[0\] _04000_ _04001_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_228_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_243_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_35_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07544_ _02764_ _03189_ _03190_ _02578_ _03191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_81_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_165_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_179_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07475_ _02597_ soc.spi_video_ram_1.write_fifo.fifo_mem\[30\]\[12\] _03122_ _02904_
+ _03123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_14_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09214_ soc.spi_video_ram_1.fifo_in_data\[11\] _04346_ _04353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_195_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06426_ _02239_ _00080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_52_1745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09145_ soc.spi_video_ram_1.state_counter\[8\] _04306_ _04308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_06357_ _02147_ soc.spi_video_ram_1.write_fifo.fifo_mem\[17\]\[13\] _02193_ _02197_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_108_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09076_ _02233_ soc.spi_video_ram_1.write_fifo.fifo_mem\[20\]\[8\] _04259_ _04268_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06288_ _02153_ soc.spi_video_ram_1.write_fifo.fifo_mem\[18\]\[16\] _02141_ _02154_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_107_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_194_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08027_ _03658_ _03660_ _03662_ _03664_ _02710_ _03665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_11_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5004 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_89_wb_clk_i clknet_5_10_0_wb_clk_i clknet_leaf_89_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_103_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5015 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5026 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09978_ soc.ram_encoder_0.input_buffer\[10\] _04869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_137_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5037 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_89_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5048 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_18_wb_clk_i clknet_5_2_0_wb_clk_i clknet_leaf_18_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_5059 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08929_ _04185_ _00636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_4325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_79_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11940_ _00999_ clknet_leaf_160_wb_clk_i soc.ram_encoder_0.input_buffer\[6\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_85_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2901 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2912 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2923 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11871_ _00930_ clknet_leaf_165_wb_clk_i net59 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_55_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2934 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_205_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2945 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_169_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2956 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10822_ soc.spi_video_ram_1.fifo_in_data\[15\] _05393_ _05397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_2967 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_232_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2978 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2989 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10753_ _04047_ _05359_ _05360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_201_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10684_ _02237_ soc.spi_video_ram_1.write_fifo.fifo_mem\[29\]\[10\] _05321_ _05322_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_205_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_220_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11305_ _00371_ clknet_leaf_196_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[26\]\[2\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_181_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12285_ _01313_ clknet_leaf_250_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[7\]\[9\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_135_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_5_20_0_wb_clk_i clknet_4_10_0_wb_clk_i clknet_5_20_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_84_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11236_ _00302_ clknet_leaf_192_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[10\]\[7\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_107_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_218_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_136_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11167_ _00233_ clknet_leaf_56_wb_clk_i soc.spi_video_ram_1.output_buffer\[23\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_6261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_171_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_231_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10118_ _04952_ _04964_ _01046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_6294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_212_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_209_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_11098_ _00164_ clknet_leaf_205_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[12\]\[7\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_5571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_114_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_236_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10049_ _04910_ _01032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_4870 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4881 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4892 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_229_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05590_ _01473_ _01489_ _01498_ _01499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_50_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07260_ _02570_ _02909_ _02910_ _02911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_84_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_108_1278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06211_ soc.spi_video_ram_1.output_buffer\[19\] soc.spi_video_ram_1.output_buffer\[16\]
+ soc.spi_video_ram_1.output_buffer\[17\] soc.spi_video_ram_1.output_buffer\[18\]
+ _01501_ _01469_ _02097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_07191_ _02629_ _02844_ _02677_ _02845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_121_1412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_30_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_185_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06142_ _02034_ soc.video_generator_1.v_count\[3\] _01861_ _02035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_145_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06073_ _01849_ _01964_ _01965_ _01966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_145_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_236_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09901_ _04812_ _02525_ _04813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_160_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09832_ soc.cpu.instruction\[3\] _04740_ _04759_ _04760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_141_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_246_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09763_ _04711_ _00945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06975_ _02612_ _02635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_6_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08714_ _03368_ _04046_ _04068_ _00538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_73_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_210_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05926_ _01594_ _01819_ _01820_ soc.cpu.PC.in\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_210_1749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09694_ soc.cpu.PC.REG.data\[10\] _04664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_67_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08645_ _04027_ _00510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_76_1509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_187_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05857_ _01722_ _01744_ _01755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_242_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_214_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_08576_ _02165_ soc.spi_video_ram_1.write_fifo.fifo_mem\[2\]\[22\] _03966_ _03991_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_82_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05788_ _01678_ _01677_ _01690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XPHY_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_126_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07527_ soc.spi_video_ram_1.write_fifo.fifo_mem\[7\]\[26\] _03175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_74_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_126_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_136_wb_clk_i clknet_5_24_0_wb_clk_i clknet_leaf_136_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_208_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07458_ _01939_ _01930_ _03106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_167_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06409_ soc.spi_video_ram_1.write_fifo.fifo_mem\[16\]\[5\] _02227_ _02217_ _02228_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_136_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_202_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_194_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07389_ _03034_ _03035_ _03037_ _02976_ _02642_ _03038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_109_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09128_ soc.spi_video_ram_1.state_counter\[1\] soc.spi_video_ram_1.state_counter\[0\]
+ soc.spi_video_ram_1.state_counter\[2\] _04297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_100_1518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_198_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_68_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_163_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09059_ _04258_ _04259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_85_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12070_ _01113_ clknet_leaf_109_wb_clk_i soc.rom_loader.current_address\[10\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_1_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11021_ _00087_ clknet_leaf_80_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[16\]\[17\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_235_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_238_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4100 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4111 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_213_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4122 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4133 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_218_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4144 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4155 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4166 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_245_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4177 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11923_ _00982_ clknet_leaf_97_wb_clk_i soc.rom_encoder_0.current_state\[1\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_4188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2720 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_166_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2731 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2742 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2753 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11854_ _00913_ clknet_leaf_96_wb_clk_i soc.rom_encoder_0.request_data_out\[15\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_32_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2764 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_233_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2775 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_226_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2786 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10805_ _02233_ soc.spi_video_ram_1.write_fifo.fifo_mem\[7\]\[8\] _05378_ _05387_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_2797 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_242_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_198_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11785_ _00846_ clknet_leaf_98_wb_clk_i soc.rom_encoder_0.output_buffer\[16\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_148_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10736_ soc.spi_video_ram_1.write_fifo.fifo_mem\[31\]\[5\] soc.spi_video_ram_1.fifo_in_data\[5\]
+ _05344_ _05350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_174_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10667_ _02221_ soc.spi_video_ram_1.write_fifo.fifo_mem\[29\]\[2\] _05310_ _05313_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_10598_ _05274_ _05268_ _05275_ _01216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_126_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12337_ _01365_ clknet_leaf_26_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[8\]\[16\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_142_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12268_ _01296_ clknet_leaf_291_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[31\]\[21\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_64_1435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11219_ _00285_ clknet_leaf_81_wb_clk_i soc.display_clks_before_active\[0\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_190_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12199_ _01227_ clknet_leaf_20_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[19\]\[10\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_96_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_6080 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6091 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_7_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_237_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06760_ soc.rom_encoder_0.output_bits_left\[3\] _02439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_5390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_23_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05711_ _01557_ _01616_ _01617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_06691_ _02396_ _00188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_224_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_188_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08430_ soc.spi_video_ram_1.write_fifo.fifo_mem\[27\]\[12\] _02242_ _03910_ _03913_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_58_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05642_ _01514_ _01515_ _01550_ _01428_ _01551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_145_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08361_ soc.spi_video_ram_1.write_fifo.fifo_mem\[26\]\[9\] _02409_ _03866_ _03876_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_05573_ _01481_ _01482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_127_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_220_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07312_ _02703_ soc.spi_video_ram_1.write_fifo.fifo_mem\[31\]\[10\] _02962_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_225_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08292_ _03838_ _00346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_149_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07243_ _02576_ _02894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_176_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_203_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07174_ soc.spi_video_ram_1.write_fifo.fifo_mem\[24\]\[6\] soc.spi_video_ram_1.write_fifo.fifo_mem\[25\]\[6\]
+ soc.spi_video_ram_1.write_fifo.fifo_mem\[26\]\[6\] soc.spi_video_ram_1.write_fifo.fifo_mem\[27\]\[6\]
+ _02763_ _02827_ _02828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_118_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_192_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_199_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06125_ _01977_ _01924_ _02005_ _02018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_69_1357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_1327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06056_ soc.video_generator_1.h_count\[8\] soc.video_generator_1.h_count\[9\] _01948_
+ _01949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_133_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_101_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_232_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09815_ _04741_ _04744_ _04745_ _04746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_115_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09746_ _04702_ _00937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_246_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06958_ _02596_ _02617_ _02618_ _02619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_100_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_227_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_223_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05909_ _01594_ _01803_ _01804_ soc.cpu.PC.in\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_2005 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09677_ soc.cpu.PC.REG.data\[5\] soc.rom_loader.current_address\[5\] _04638_ _04652_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_27_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_317_wb_clk_i clknet_5_0_0_wb_clk_i clknet_leaf_317_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_2016 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06889_ _02553_ _02554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_43_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2027 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2038 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_243_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2049 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08628_ _02155_ soc.spi_video_ram_1.write_fifo.fifo_mem\[30\]\[17\] _04011_ _04019_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_215_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_93_1631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_199_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08559_ _03982_ _00469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_243_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_196_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11570_ _00636_ clknet_leaf_248_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[22\]\[6\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_180_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_210_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_168_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10521_ _01565_ _05228_ _05230_ _01184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_122_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xcaravel_hack_soc_201 wbs_dat_o[9] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_10452_ soc.cpu.PC.REG.data\[0\] soc.cpu.PC.REG.data\[1\] _05177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_52_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_1424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xcaravel_hack_soc_212 wbs_dat_o[20] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xcaravel_hack_soc_223 wbs_dat_o[31] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_136_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_201_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_182_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_174_1405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_30_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10383_ _02233_ soc.spi_video_ram_1.write_fifo.fifo_mem\[6\]\[8\] _05124_ _05133_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_178_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12122_ _01150_ clknet_leaf_317_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[6\]\[14\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_leaf_33_wb_clk_i clknet_5_9_0_wb_clk_i clknet_leaf_33_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_124_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_12053_ net31 clknet_leaf_87_wb_clk_i soc.rom_encoder_0.data_out\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_151_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11004_ _00070_ clknet_leaf_222_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[16\]\[0\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_81_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_219_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_206_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_209_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11906_ _00965_ clknet_leaf_124_wb_clk_i soc.cpu.DMuxJMP.sel\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_61_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11837_ _00896_ clknet_leaf_123_wb_clk_i soc.rom_encoder_0.input_buffer\[11\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_199_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_187_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1860 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1871 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_202_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_183_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1882 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1893 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11768_ _00829_ clknet_leaf_69_wb_clk_i soc.spi_video_ram_1.sram_sck_fall_edge vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_109_1384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_187_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_186_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_159_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10719_ _03160_ _05324_ _05340_ _01272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_201_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11699_ _00760_ clknet_5_22_0_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[9\]\[1\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_228_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_155_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_196_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_170_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07930_ _01898_ _02625_ _03572_ _02734_ _03573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_116_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_233_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07861_ _02700_ _03504_ _03505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_110_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_111_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09600_ soc.rom_encoder_0.input_buffer\[3\] _04586_ _04601_ _04602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_84_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06812_ soc.ram_encoder_0.request_write _02483_ _02487_ _02488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_110_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07792_ _02984_ _03433_ _03436_ _03437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_209_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09531_ _01380_ _04553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_42_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06743_ _02427_ _00209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_3_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_225_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_184_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09462_ _04473_ _04507_ _04508_ _00847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06674_ _02173_ soc.spi_video_ram_1.write_fifo.fifo_mem\[12\]\[26\] _02356_ _02385_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_129_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08413_ soc.spi_video_ram_1.write_fifo.fifo_mem\[27\]\[4\] _02399_ _03899_ _03904_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_149_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05625_ soc.spi_video_ram_1.output_buffer\[20\] _01534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09393_ _04455_ _00831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08344_ _03867_ _00369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05556_ soc.spi_video_ram_1.buffer_index\[4\] _01464_ _01465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_240_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_193_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08275_ _02558_ _03827_ _03828_ _00339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_138_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05487_ _01399_ _01401_ _01402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_123_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07226_ _02650_ _02877_ _02618_ _02878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_138_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_193_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_175_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xclkbuf_4_1_0_wb_clk_i clknet_3_0_0_wb_clk_i clknet_4_1_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_69_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07157_ _02596_ _02811_ _02812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_121_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_238_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06108_ _01977_ _02000_ _01978_ _01922_ _02001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_175_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07088_ _02744_ soc.spi_video_ram_1.write_fifo.fifo_mem\[6\]\[3\] _02745_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_82_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06039_ _01930_ _01931_ _01859_ _01932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_105_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_236_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09729_ net60 _04677_ _04692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_leaf_151_wb_clk_i clknet_5_30_0_wb_clk_i clknet_leaf_151_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_90_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_242_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11622_ _00688_ clknet_leaf_47_wb_clk_i _00000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_106_1502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_11_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_230_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_211_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_168_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11553_ _00619_ clknet_leaf_23_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[25\]\[18\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_184_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10504_ soc.cpu.PC.in\[14\] _05188_ _05201_ _05217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_52_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_144_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11484_ _00550_ clknet_leaf_185_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[24\]\[7\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_170_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10435_ _01699_ _01736_ _05161_ _05162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_109_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_178_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10366_ _05123_ _05124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_48_1249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12105_ _01133_ net85 soc.cpu.ALU.x\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_174_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_139_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10297_ soc.rom_loader.current_address\[5\] _05080_ _05082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_156_1680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_97_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12036_ _01095_ clknet_leaf_302_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[5\]\[24\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_leaf_239_wb_clk_i clknet_5_16_0_wb_clk_i clknet_leaf_239_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_61_1438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_77_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_238_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_168_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_207_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3070 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3081 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_234_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3092 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_146_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_18_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06390_ soc.spi_video_ram_1.write_fifo.write_pointer\[1\] _01405_ _02214_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_226_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_175_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_193_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_187_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_159_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_204_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08060_ soc.spi_video_ram_1.write_fifo.fifo_mem\[11\]\[8\] _02407_ _03680_ _03689_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_198_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07011_ soc.spi_video_ram_1.output_buffer\[21\] _02670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_179_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_179_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08962_ _04202_ _00652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_192_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_237_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07913_ _02689_ soc.spi_video_ram_1.write_fifo.fifo_mem\[22\]\[21\] _03555_ _02593_
+ _03556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_97_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_25_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08893_ _04165_ _00620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_151_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_131_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07844_ _02984_ _03484_ _03487_ _03488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_56_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07775_ _02907_ _03419_ _03420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_72_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_83_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09514_ _02268_ soc.cpu.AReg.data\[9\] _01459_ _04542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_25_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06726_ soc.spi_video_ram_1.write_fifo.fifo_mem\[14\]\[15\] _02248_ _02412_ _02419_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_37_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_224_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09445_ soc.rom_encoder_0.output_buffer\[14\] _04479_ _04495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06657_ _02376_ _00174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_129_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_244_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_05608_ soc.spi_video_ram_1.output_buffer\[8\] soc.spi_video_ram_1.output_buffer\[9\]
+ _01468_ _01517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_240_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_185_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09376_ soc.spi_video_ram_1.state_sram_clk_counter\[6\] _04443_ _04445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_36_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06588_ soc.spi_video_ram_1.fifo_in_address\[1\] _02337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_212_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08327_ _03856_ _00363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_16_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05539_ _01403_ soc.spi_video_ram_1.write_fifo.write_pointer\[2\] _01445_ _01449_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_197_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08258_ soc.ram_encoder_0.output_buffer\[12\] _03814_ _03815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07209_ soc.spi_video_ram_1.write_fifo.fifo_mem\[8\]\[8\] soc.spi_video_ram_1.write_fifo.fifo_mem\[9\]\[8\]
+ soc.spi_video_ram_1.write_fifo.fifo_mem\[10\]\[8\] soc.spi_video_ram_1.write_fifo.fifo_mem\[11\]\[8\]
+ _02575_ _02578_ _02861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_152_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08189_ _03760_ _00321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_88_1574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10220_ _02229_ soc.spi_video_ram_1.write_fifo.fifo_mem\[5\]\[6\] _05030_ _05037_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_3_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10151_ _04986_ _04988_ _04989_ _01054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_171_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5901 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5912 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5923 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_47_1282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10082_ net2 _04834_ _04936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_134_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5934 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5945 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_199_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_48_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5956 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_216_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5967 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5978 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_87_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5989 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_1501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_210_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_244_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10984_ _00050_ clknet_leaf_248_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[17\]\[9\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_216_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_243_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11605_ _00671_ clknet_leaf_306_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[21\]\[12\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_169_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_184_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11536_ _00602_ clknet_leaf_180_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[25\]\[1\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_157_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_221_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_172_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_171_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11467_ _00533_ clknet_leaf_29_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[15\]\[19\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_99_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10418_ _02268_ soc.spi_video_ram_1.write_fifo.fifo_mem\[6\]\[25\] _05123_ _05151_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_11398_ _00464_ clknet_leaf_220_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[2\]\[8\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_180_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10349_ _01736_ _05103_ _05114_ _01128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_124_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_193_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_234_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_117_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12019_ _01078_ clknet_leaf_243_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[5\]\[7\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_239_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05890_ _01782_ _01785_ _01786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_94_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_187_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07560_ _02586_ _03192_ _03197_ _03206_ _03207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_34_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_235_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06511_ _02293_ _00111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_206_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07491_ _02679_ _03139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_61_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09230_ _04362_ _00760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_94_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06442_ soc.spi_video_ram_1.fifo_in_address\[0\] _02250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_222_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_167_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09161_ soc.video_generator_1.v_count\[1\] _04313_ _04320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06373_ _02163_ soc.spi_video_ram_1.write_fifo.fifo_mem\[17\]\[21\] _02181_ _02205_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_72_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08112_ soc.video_generator_1.h_count\[3\] soc.video_generator_1.h_count\[2\] _03715_
+ _03717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_33_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09092_ _04276_ _00708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_222_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08043_ _03679_ _03680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_102_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_147_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_190_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_198_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_200_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_150_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09994_ soc.ram_encoder_0.request_data_out\[0\] soc.ram_encoder_0.data_out\[0\] _04880_
+ _04882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_157_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_213_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08945_ soc.spi_video_ram_1.write_fifo.fifo_mem\[22\]\[14\] _04052_ _04189_ _04194_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_135_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_213_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08876_ soc.spi_video_ram_1.write_fifo.fifo_mem\[25\]\[11\] _02414_ _04155_ _04157_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_97_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3806 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3817 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_229_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3828 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07827_ _02918_ _03448_ _03471_ _03472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_85_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3839 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_229_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_178_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_245_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_246_1501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_226_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_211_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07758_ _03021_ soc.spi_video_ram_1.write_fifo.fifo_mem\[13\]\[15\] _03402_ _03024_
+ _03403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_77_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_231_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_53_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06709_ _02408_ _00194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_225_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07689_ soc.spi_video_ram_1.write_fifo.fifo_mem\[23\]\[24\] _03335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_1571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09428_ soc.rom_encoder_0.request_address\[9\] _02520_ _04460_ soc.rom_encoder_0.output_buffer\[6\]
+ _04481_ _04482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_0_1593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_241_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_198_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09359_ soc.spi_video_ram_1.state_sram_clk_counter\[0\] _04431_ _04433_ _04434_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_60_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_240_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11321_ _00387_ clknet_leaf_23_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[26\]\[18\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_177_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_153_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_5_10_0_wb_clk_i clknet_4_5_0_wb_clk_i clknet_5_10_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_11252_ _00318_ clknet_leaf_237_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[10\]\[23\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_181_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10203_ soc.hack_clock_0.counter\[5\] _05024_ _05027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_162_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_106_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11183_ _00249_ clknet_leaf_59_wb_clk_i soc.spi_video_ram_1.output_buffer\[7\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_6421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_238_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10134_ _04952_ _04976_ _01050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_7_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_122_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5720 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_122_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5731 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5742 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5753 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10065_ _04919_ _04921_ soc.ram_encoder_0.initializing_step\[0\] _04922_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_7_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5764 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_1702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_5775 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5786 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_235_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_5797 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_188_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_169_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_217_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_1410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_229_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_182_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10967_ _00033_ clknet_leaf_241_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[18\]\[21\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_56_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_204_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_206_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10898_ _05437_ _01354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_31_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_200_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_11519_ _00585_ clknet_leaf_39_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[23\]\[13\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_116_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_236_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_254_wb_clk_i clknet_5_7_0_wb_clk_i clknet_leaf_254_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_125_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_153_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_125_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_217_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06991_ _02612_ _02651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_113_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08730_ _04078_ _00544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05942_ _01594_ _01834_ _01835_ soc.cpu.PC.in\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08661_ _04036_ _00517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_230_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05873_ _01670_ soc.cpu.ALU.x\[11\] _01770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_67_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07612_ soc.spi_video_ram_1.write_fifo.fifo_mem\[7\]\[25\] _03259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_208_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08592_ _03999_ _04000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_82_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_241_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_198_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07543_ _02591_ soc.spi_video_ram_1.write_fifo.fifo_mem\[20\]\[13\] _03190_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_207_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_210_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_201_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07474_ _02931_ _03121_ _03122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_223_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09213_ _04341_ _01767_ _04352_ _00753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_194_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06425_ soc.spi_video_ram_1.write_fifo.fifo_mem\[16\]\[10\] _02237_ _02238_ _02239_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_33_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09144_ _04294_ _04306_ _04307_ _00729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_241_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06356_ _02196_ _00053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_163_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09075_ _04267_ _00700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_135_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06287_ soc.spi_video_ram_1.fifo_in_address\[0\] _02153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_190_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08026_ _02685_ _03663_ _03579_ _03664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_146_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_163_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_235_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5005 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5016 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_104_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09977_ _04867_ _04848_ _04868_ _01002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_131_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5027 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5038 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5049 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_118_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08928_ soc.spi_video_ram_1.write_fifo.fifo_mem\[22\]\[6\] _02403_ _04178_ _04185_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_4326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_217_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08859_ soc.spi_video_ram_1.write_fifo.fifo_mem\[25\]\[3\] _02397_ _04144_ _04148_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_3625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2902 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_233_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2913 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11870_ _00929_ clknet_leaf_165_wb_clk_i net58 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_leaf_58_wb_clk_i clknet_5_12_0_wb_clk_i clknet_leaf_58_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_3658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2924 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2935 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2946 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10821_ _03323_ _05392_ _05396_ _01318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_2957 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_60_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2968 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2979 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_41_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10752_ _05343_ _05359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_197_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_207_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_200_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_186_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_231_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10683_ _05309_ _05321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_125_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_199_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_127_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11304_ _00370_ clknet_leaf_187_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[26\]\[1\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12284_ _01312_ clknet_leaf_244_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[7\]\[8\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_4_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11235_ _00301_ clknet_leaf_203_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[10\]\[6\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_136_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_214_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11166_ _00232_ clknet_leaf_149_wb_clk_i soc.ram_encoder_0.output_buffer\[1\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_84_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_95_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10117_ soc.ram_data_out\[8\] _04927_ _04963_ _04964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_6284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_49_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_4_14_0_wb_clk_i clknet_3_7_0_wb_clk_i clknet_4_14_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XTAP_6295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11097_ _00163_ clknet_leaf_203_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[12\]\[6\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_5561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10048_ soc.ram_encoder_0.request_address\[10\] soc.ram_encoder_0.address\[10\] _04900_
+ _04910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_3_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_231_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4860 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4871 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4882 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4893 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_236_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_223_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11999_ _01058_ clknet_leaf_164_wb_clk_i soc.ram_encoder_0.current_state\[2\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_91_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_225_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_205_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_182_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_182_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06210_ _02089_ _02091_ _02095_ _02096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_34_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_192_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07190_ _02606_ _02833_ _02843_ _02844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_77_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06141_ soc.video_generator_1.v_count\[4\] _02034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_117_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_172_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06072_ _01939_ _01940_ _01932_ _01965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_104_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09900_ _02436_ _02454_ _04812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_99_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_119_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09831_ _04741_ _04757_ _04758_ _04759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_154_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_236_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09762_ _02242_ soc.spi_video_ram_1.write_fifo.fifo_mem\[3\]\[12\] _04708_ _04711_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06974_ _02634_ _00233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_80_1485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05925_ _01552_ soc.cpu.instruction\[13\] soc.cpu.AReg.data\[13\] _01591_ _01820_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_08713_ _04067_ _04048_ _04068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09693_ _04663_ _00923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_66_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_215_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08644_ _02171_ soc.spi_video_ram_1.write_fifo.fifo_mem\[30\]\[25\] _03999_ _04027_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_2209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05856_ _01732_ _01733_ _01729_ _01746_ _01754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XPHY_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_199_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08575_ _03990_ _00477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05787_ _01684_ _01688_ _01689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XPHY_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_165_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_74_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_165_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07526_ soc.spi_video_ram_1.write_fifo.fifo_mem\[0\]\[26\] soc.spi_video_ram_1.write_fifo.fifo_mem\[1\]\[26\]
+ soc.spi_video_ram_1.write_fifo.fifo_mem\[2\]\[26\] soc.spi_video_ram_1.write_fifo.fifo_mem\[3\]\[26\]
+ _02919_ _02577_ _03174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_211_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_161_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07457_ _03015_ _03104_ _03105_ _00244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_50_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06408_ soc.spi_video_ram_1.fifo_in_data\[5\] _02227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_07388_ _02696_ soc.spi_video_ram_1.write_fifo.fifo_mem\[28\]\[11\] _03036_ _03037_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xclkbuf_leaf_176_wb_clk_i clknet_5_23_0_wb_clk_i clknet_leaf_176_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_109_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_176_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09127_ soc.spi_video_ram_1.state_counter\[1\] soc.spi_video_ram_1.state_counter\[0\]
+ soc.spi_video_ram_1.state_counter\[2\] _04296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_210_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06339_ _02187_ _00045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xclkbuf_leaf_105_wb_clk_i clknet_5_14_0_wb_clk_i clknet_leaf_105_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_178_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_191_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_194_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09058_ _04257_ _04258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_68_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08009_ soc.spi_video_ram_1.write_fifo.fifo_mem\[28\]\[17\] soc.spi_video_ram_1.write_fifo.fifo_mem\[29\]\[17\]
+ soc.spi_video_ram_1.write_fifo.fifo_mem\[30\]\[17\] soc.spi_video_ram_1.write_fifo.fifo_mem\[31\]\[17\]
+ _02726_ _03041_ _03648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_123_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_2_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_150_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11020_ _00086_ clknet_leaf_75_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[16\]\[16\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_215_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_1317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4101 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4112 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4123 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4134 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4145 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4156 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_4167 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4178 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11922_ _00981_ clknet_leaf_97_wb_clk_i soc.rom_encoder_0.current_state\[0\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_4189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2710 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_218_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2721 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_205_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_185_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2732 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2743 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11853_ _00912_ clknet_leaf_100_wb_clk_i soc.rom_encoder_0.request_data_out\[14\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2754 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2765 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2776 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2787 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10804_ _05386_ _01311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_11784_ _00845_ clknet_leaf_102_wb_clk_i soc.rom_encoder_0.output_buffer\[15\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2798 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_226_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_201_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10735_ _05349_ _01279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_14_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_220_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_174_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10666_ _05312_ _01247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_167_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_127_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10597_ soc.gpio_i_stored\[3\] _05268_ _02053_ _05275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_12_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12336_ _01364_ clknet_leaf_9_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[8\]\[15\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_127_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_181_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12267_ _01295_ clknet_leaf_56_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[31\]\[20\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_218_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_233_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11218_ _00284_ clknet_leaf_269_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[11\]\[28\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_9_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_12198_ _01226_ clknet_leaf_256_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[19\]\[9\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xoutput80 net80 io_out[37] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_96_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11149_ _00215_ clknet_leaf_125_wb_clk_i net65 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_228_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6070 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6081 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6092 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_49_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_5_3_0_wb_clk_i clknet_4_1_0_wb_clk_i clknet_5_3_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_05710_ _01558_ soc.cpu.ALU.x\[2\] _01616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06690_ soc.spi_video_ram_1.write_fifo.fifo_mem\[14\]\[2\] _02395_ _02391_ _02396_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_110_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05641_ soc.spi_video_ram_1.buffer_index\[4\] _01527_ _01549_ _01463_ _01550_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_36_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08360_ _03875_ _00377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05572_ _01476_ _01479_ _01480_ _01467_ _01481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
Xclkbuf_leaf_3_wb_clk_i clknet_5_2_0_wb_clk_i clknet_leaf_3_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_07311_ soc.spi_video_ram_1.write_fifo.fifo_mem\[24\]\[10\] soc.spi_video_ram_1.write_fifo.fifo_mem\[25\]\[10\]
+ soc.spi_video_ram_1.write_fifo.fifo_mem\[26\]\[10\] soc.spi_video_ram_1.write_fifo.fifo_mem\[27\]\[10\]
+ _02574_ _02592_ _02961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_60_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08291_ _02132_ soc.spi_video_ram_1.write_fifo.fifo_mem\[1\]\[6\] _03831_ _03838_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_127_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07242_ _02679_ _02893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_20_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_242_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07173_ _02646_ _02827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_121_1243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06124_ _01977_ _01924_ _02017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_195_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06055_ soc.video_generator_1.h_count\[8\] _01837_ _01948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_132_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09814_ net5 _04566_ _04745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_115_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_246_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09745_ _02225_ soc.spi_video_ram_1.write_fifo.fifo_mem\[3\]\[4\] _04697_ _04702_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_210_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06957_ _02601_ _02618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_86_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05908_ _01552_ _01598_ soc.cpu.AReg.data\[12\] _01591_ _01804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XTAP_2006 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09676_ _04651_ _00918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06888_ soc.ram_encoder_0.toggled_sram_sck _02489_ _02498_ _02552_ _02553_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__nand4_1
XTAP_2017 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2028 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_242_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2039 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05839_ _01732_ _01733_ _01729_ _01738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08627_ _04018_ _00501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_110_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_19_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_230_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08558_ _02147_ soc.spi_video_ram_1.write_fifo.fifo_mem\[2\]\[13\] _03978_ _03982_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_74_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_208_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07509_ soc.spi_video_ram_1.write_fifo.fifo_mem\[31\]\[26\] _03157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_08489_ _03932_ _03945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_51_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10520_ soc.ram_encoder_0.address\[1\] _05228_ _05230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_161_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_156_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_221_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_202_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10451_ _05171_ _05175_ _05176_ _01167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xcaravel_hack_soc_202 wbs_dat_o[10] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_136_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xcaravel_hack_soc_213 wbs_dat_o[21] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_136_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xcaravel_hack_soc_224 io_oeb[26] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_163_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10382_ _05132_ _01143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_184_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12121_ _01149_ clknet_leaf_314_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[6\]\[13\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_237_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_219_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_151_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12052_ net30 clknet_leaf_112_wb_clk_i soc.rom_encoder_0.data_out\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_151_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_78_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_238_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11003_ _00069_ clknet_leaf_278_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[17\]\[28\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_46_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_73_wb_clk_i clknet_5_8_0_wb_clk_i clknet_leaf_73_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_120_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_237_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_111_1412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_234_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11905_ _00964_ clknet_leaf_127_wb_clk_i soc.cpu.DMuxJMP.sel\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_46_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_185_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_233_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_226_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11836_ _00895_ clknet_leaf_125_wb_clk_i soc.rom_encoder_0.input_buffer\[10\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1850 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1861 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_42_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1872 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1894 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11767_ _00828_ clknet_leaf_63_wb_clk_i soc.spi_video_ram_1.sram_sck_rise_edge vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
X_10718_ soc.spi_video_ram_1.fifo_in_address\[10\] _05325_ _05340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_11698_ _00759_ clknet_leaf_191_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[9\]\[0\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_179_1317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10649_ soc.spi_video_ram_1.write_fifo.fifo_mem\[19\]\[23\] _04065_ _05277_ _05303_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_127_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_200_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_192_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_12319_ _01347_ clknet_leaf_115_wb_clk_i soc.ram_encoder_0.data_out\[14\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_142_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_244_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_190_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07860_ soc.spi_video_ram_1.write_fifo.fifo_mem\[5\]\[22\] _03504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_229_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06811_ _02484_ _02486_ _02487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_151_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07791_ _02689_ soc.spi_video_ram_1.write_fifo.fifo_mem\[20\]\[23\] _03435_ _02742_
+ _03436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_49_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06742_ soc.spi_video_ram_1.write_fifo.fifo_mem\[14\]\[23\] _02264_ _02390_ _02427_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_09530_ soc.spi_video_ram_1.fifo_read_request _04551_ soc.spi_video_ram_1.fifo_write_request
+ _04552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_224_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_188_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09461_ soc.rom_encoder_0.output_buffer\[17\] _04479_ _04508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_58_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_06673_ _02384_ _00182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_97_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05624_ _01501_ _01508_ _01532_ _01533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_08412_ _03903_ _00401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_212_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09392_ net9 soc.spi_video_ram_1.read_value\[0\] _04454_ _04455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_75_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08343_ soc.spi_video_ram_1.write_fifo.fifo_mem\[26\]\[0\] _02310_ _03866_ _03867_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_05555_ soc.spi_video_ram_1.buffer_index\[2\] _01463_ _01464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_33_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_225_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_149_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_1485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08274_ soc.ram_encoder_0.output_buffer\[19\] _02555_ _03828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_138_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05486_ soc.spi_video_ram_1.write_fifo.read_pointer\[1\] _01400_ _01401_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_203_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07225_ soc.spi_video_ram_1.write_fifo.fifo_mem\[20\]\[8\] soc.spi_video_ram_1.write_fifo.fifo_mem\[21\]\[8\]
+ soc.spi_video_ram_1.write_fifo.fifo_mem\[22\]\[8\] soc.spi_video_ram_1.write_fifo.fifo_mem\[23\]\[8\]
+ _02591_ _02593_ _02877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_118_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_140_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_192_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07156_ soc.spi_video_ram_1.write_fifo.fifo_mem\[28\]\[5\] soc.spi_video_ram_1.write_fifo.fifo_mem\[29\]\[5\]
+ soc.spi_video_ram_1.write_fifo.fifo_mem\[30\]\[5\] soc.spi_video_ram_1.write_fifo.fifo_mem\[31\]\[5\]
+ _02635_ _02636_ _02811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_145_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06107_ _01986_ _01988_ _01999_ _01967_ _02000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_07087_ _02590_ _02744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_161_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06038_ soc.video_generator_1.v_count\[3\] _01931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_216_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_232_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_219_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07989_ _03577_ _03628_ _02720_ _03629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_216_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09728_ soc.ram_encoder_0.output_buffer\[18\] _03814_ _03788_ soc.ram_encoder_0.request_data_out\[14\]
+ _03817_ _04691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_41_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_243_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09659_ _04638_ _04639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_16_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_215_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_16_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_188_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_191_wb_clk_i clknet_5_22_0_wb_clk_i clknet_leaf_191_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_231_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_1451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_243_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11621_ _00687_ clknet_leaf_274_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[21\]\[28\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_54_1424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_196_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_223_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_180_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11552_ _00618_ clknet_leaf_22_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[25\]\[17\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_184_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_156_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_195_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10503_ soc.cpu.PC.REG.data\[14\] _05215_ _05216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_11483_ _00549_ clknet_leaf_201_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[24\]\[6\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_137_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10434_ _01666_ _01680_ _01713_ _05160_ _05161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_152_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10365_ _05122_ _05123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_124_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_124_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12104_ _01132_ net85 soc.cpu.ALU.x\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10296_ soc.rom_loader.current_address\[5\] _05080_ _05081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_124_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_156_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_191_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_239_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_12035_ _01094_ clknet_leaf_287_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[5\]\[23\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_2_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_215_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_20_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_279_wb_clk_i clknet_5_4_0_wb_clk_i clknet_leaf_279_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_206_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_189_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3060 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_208_wb_clk_i clknet_5_22_0_wb_clk_i clknet_leaf_208_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_3071 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3082 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3093 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_146_1327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_181_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_221_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11819_ _00878_ clknet_leaf_71_wb_clk_i soc.spi_video_ram_1.write_fifo.read_pointer\[1\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_222_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_186_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_179_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07010_ _02669_ _00234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_127_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_196_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_183_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08961_ soc.spi_video_ram_1.write_fifo.fifo_mem\[22\]\[22\] _04063_ _04177_ _04202_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_29_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07912_ _02651_ _03554_ _03555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_64_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_233_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08892_ soc.spi_video_ram_1.write_fifo.fifo_mem\[25\]\[19\] _02341_ _04155_ _04165_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_25_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07843_ _02764_ soc.spi_video_ram_1.write_fifo.fifo_mem\[20\]\[22\] _03486_ _02742_
+ _03487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_97_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_245_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07774_ soc.spi_video_ram_1.write_fifo.fifo_mem\[5\]\[15\] _03419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_42_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09513_ _04541_ _00865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_225_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06725_ _02418_ _00200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_52_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_20_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09444_ soc.rom_encoder_0.request_address\[13\] _02520_ _04460_ soc.rom_encoder_0.output_buffer\[10\]
+ _04493_ _04494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_06656_ _02155_ soc.spi_video_ram_1.write_fifo.fifo_mem\[12\]\[17\] _02368_ _02376_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_168_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_213_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_05607_ _01469_ _01470_ _01516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_06587_ _02336_ _00144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09375_ _04443_ _04444_ _00823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_240_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08326_ _02167_ soc.spi_video_ram_1.write_fifo.fifo_mem\[1\]\[23\] _03830_ _03856_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_05538_ _01398_ _01441_ _01447_ _01448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_162_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08257_ _02480_ _02498_ _03779_ _03814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_21_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05469_ _01382_ _01383_ _01384_ _01385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_166_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_193_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07208_ _01510_ _02676_ _02848_ _02860_ _00240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_101_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08188_ _02173_ soc.spi_video_ram_1.write_fifo.fifo_mem\[10\]\[26\] _03731_ _03760_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_88_1542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_119_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07139_ _02685_ _02794_ _02720_ _02795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_238_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10150_ net81 _04986_ _01395_ _04989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_121_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5902 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5913 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10081_ soc.ram_encoder_0.request_data_out\[1\] _04930_ _04935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_88_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5924 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_173_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_5935 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5946 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5957 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5968 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5979 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_75_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_301_wb_clk_i clknet_5_1_0_wb_clk_i clknet_leaf_301_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_10983_ _00049_ clknet_5_23_0_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[17\]\[8\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_95_1535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_128_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_203_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_230_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11604_ _00670_ clknet_leaf_34_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[21\]\[11\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_180_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_223_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11535_ _00601_ clknet_leaf_184_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[25\]\[0\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_8_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_184_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_156_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_139_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11466_ _00532_ clknet_leaf_22_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[15\]\[18\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_183_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10417_ _05150_ _01160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_87_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11397_ _00463_ clknet_leaf_200_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[2\]\[7\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_125_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_180_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_180_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10348_ soc.cpu.ALU.x\[8\] _05109_ _05114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10279_ soc.rom_loader.current_address\[0\] _01119_ _05069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_174_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_230_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_12018_ _01077_ clknet_leaf_246_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[5\]\[6\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_79_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_238_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_207_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_234_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06510_ _02145_ soc.spi_video_ram_1.write_fifo.fifo_mem\[0\]\[12\] _02290_ _02293_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_146_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07490_ _02712_ soc.spi_video_ram_1.write_fifo.fifo_mem\[12\]\[12\] _02943_ _03138_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_228_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06441_ _02249_ _00085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_146_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_146_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_226_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_241_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09160_ _04313_ _04317_ _04319_ _00733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_06372_ _02204_ _00061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_187_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08111_ _03713_ _03716_ _00287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_159_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09091_ _02248_ soc.spi_video_ram_1.write_fifo.fifo_mem\[20\]\[15\] _04270_ _04276_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_50_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08042_ _03678_ _03679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_190_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_1753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_239_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_171_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09993_ _03816_ _04880_ _04881_ _01005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_66_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_192_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_118_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08944_ _04193_ _00643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_69_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08875_ _04156_ _00611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_56_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3807 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3818 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07826_ _02656_ _03457_ _03470_ _03471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_3829 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_44_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07757_ _02919_ soc.spi_video_ram_1.write_fifo.fifo_mem\[12\]\[15\] _03402_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_84_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_71_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06708_ soc.spi_video_ram_1.write_fifo.fifo_mem\[14\]\[8\] _02407_ _02391_ _02408_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_168_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07688_ _02958_ _03330_ _03333_ _02706_ _03334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_73_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09427_ soc.rom_encoder_0.request_data_out\[2\] _03767_ _04481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_06639_ _02138_ soc.spi_video_ram_1.write_fifo.fifo_mem\[12\]\[9\] _02357_ _02367_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_240_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_212_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09358_ soc.spi_video_ram_1.current_state\[2\] net68 _04433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_139_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_1476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08309_ _03847_ _00354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09289_ _04393_ _04394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_138_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11320_ _00386_ clknet_leaf_23_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[26\]\[17\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_10_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_158_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11251_ _00317_ clknet_leaf_252_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[10\]\[22\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_107_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_162_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10202_ _05017_ _05026_ _01069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_136_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11182_ _00248_ clknet_leaf_62_wb_clk_i soc.spi_video_ram_1.output_buffer\[8\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_6400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_192_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10133_ soc.ram_data_out\[12\] _04928_ _04975_ _04976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_161_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5710 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5721 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5732 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_216_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5743 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10064_ _04830_ _04920_ _04921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_76_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_6499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5754 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5765 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5776 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_102_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5787 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5798 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_236_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_169_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_235_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_245_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_216_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_189_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10966_ _00032_ clknet_leaf_51_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[18\]\[20\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_232_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_245_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10897_ soc.spi_video_ram_1.write_fifo.fifo_mem\[8\]\[5\] soc.spi_video_ram_1.fifo_in_data\[5\]
+ _05431_ _05437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_182_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_227_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_231_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_157_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11518_ _00584_ clknet_leaf_306_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[23\]\[12\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_171_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11449_ _00515_ clknet_leaf_222_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[15\]\[1\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_113_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_193_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_119_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_234_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_294_wb_clk_i clknet_5_4_0_wb_clk_i clknet_leaf_294_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06990_ _02569_ _02650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_132_1702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05941_ _01552_ soc.cpu.instruction\[14\] soc.cpu.AReg.data\[14\] _01591_ _01835_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XTAP_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_239_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_187_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05872_ _01758_ _01761_ _01763_ _01682_ _01769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_08660_ soc.spi_video_ram_1.write_fifo.fifo_mem\[15\]\[3\] _02397_ _04032_ _04036_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_187_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07611_ _02920_ soc.spi_video_ram_1.write_fifo.fifo_mem\[4\]\[25\] _03257_ _03024_
+ _03258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_26_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08591_ _03998_ _03999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_53_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_235_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07542_ soc.spi_video_ram_1.write_fifo.fifo_mem\[21\]\[13\] _03189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_07473_ soc.spi_video_ram_1.write_fifo.fifo_mem\[31\]\[12\] _03121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_222_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_161_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09212_ soc.spi_video_ram_1.fifo_in_data\[10\] _04346_ _04352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_37_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06424_ _02215_ _02238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_210_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_124_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06355_ _02145_ soc.spi_video_ram_1.write_fifo.fifo_mem\[17\]\[12\] _02193_ _02196_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_52_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09143_ soc.spi_video_ram_1.state_counter\[7\] _04304_ _04307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_206_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09074_ _02231_ soc.spi_video_ram_1.write_fifo.fifo_mem\[20\]\[7\] _04259_ _04267_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06286_ _02152_ _00027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_147_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_198_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_163_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_159_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08025_ soc.spi_video_ram_1.write_fifo.fifo_mem\[12\]\[16\] soc.spi_video_ram_1.write_fifo.fifo_mem\[13\]\[16\]
+ soc.spi_video_ram_1.write_fifo.fifo_mem\[14\]\[16\] soc.spi_video_ram_1.write_fifo.fifo_mem\[15\]\[16\]
+ _02717_ _02682_ _03663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_200_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_116_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_190_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5006 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09976_ soc.ram_encoder_0.input_buffer\[5\] _04847_ _04248_ _04868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_5017 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_77_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5028 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_5039 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_162_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_131_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08927_ _04184_ _00635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_103_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_4305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_57_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_218_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08858_ _04147_ _00603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07809_ _02688_ _03453_ _03454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2903 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_211_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2914 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08789_ _04109_ _04110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XTAP_2925 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_217_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_1319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2936 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10820_ soc.spi_video_ram_1.fifo_in_data\[14\] _05393_ _05396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_96_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2947 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2958 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2969 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_214_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_98_wb_clk_i clknet_5_14_0_wb_clk_i clknet_leaf_98_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_10751_ _05355_ _05358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_92_1549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_241_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_198_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_183_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_213_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_27_wb_clk_i clknet_5_8_0_wb_clk_i clknet_leaf_27_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_10682_ _05320_ _01255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_90_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_224_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_187_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_9_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_224_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_107_1483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_200_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_154_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_177_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11303_ _00369_ clknet_leaf_184_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[26\]\[0\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_142_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12283_ _01311_ clknet_leaf_244_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[7\]\[7\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_84_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11234_ _00300_ clknet_leaf_205_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[10\]\[5\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_135_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_106_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11165_ _00231_ clknet_leaf_149_wb_clk_i soc.ram_encoder_0.output_buffer\[2\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_6241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_122_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_6263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_49_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10116_ _04857_ _04947_ _04948_ _04962_ _04963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_114_1410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11096_ _00162_ clknet_leaf_224_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[12\]\[5\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_6285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10047_ _04909_ _01031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_62_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_23_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4850 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4861 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4872 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_1438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_212_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4883 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_5_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4894 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_217_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11998_ _01057_ clknet_leaf_165_wb_clk_i soc.ram_encoder_0.current_state\[1\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_147_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_204_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_147_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10949_ _00015_ clknet_leaf_140_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[18\]\[3\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_147_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_242_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_143_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_203_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_125_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_203_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06140_ _01836_ soc.video_generator_1.h_count\[6\] _02032_ _02033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_129_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_184_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_219_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06071_ _01853_ _01849_ _01964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_201_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_99_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09830_ net8 _04566_ _04758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_113_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_141_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09761_ _04710_ _00944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_140_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_132_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06973_ soc.spi_video_ram_1.output_buffer\[23\] _02628_ _02633_ _02634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_39_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08712_ soc.spi_video_ram_1.fifo_in_address\[8\] _04067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_05924_ _01654_ _01818_ _01819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_09692_ _04662_ soc.rom_encoder_0.request_address\[9\] _04617_ _04663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_67_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_230_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08643_ _04026_ _00509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_6_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05855_ _01595_ _01752_ _01753_ soc.cpu.PC.in\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_54_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_94_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08574_ _02163_ soc.spi_video_ram_1.write_fifo.fifo_mem\[2\]\[21\] _03966_ _03990_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XPHY_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_05786_ _01561_ _01687_ _01688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XPHY_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_54_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_35_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07525_ _02984_ _03166_ _03172_ _02585_ _03173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_39_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_223_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_161_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_228_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_194_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07456_ soc.spi_video_ram_1.output_buffer\[12\] _02676_ _03105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_211_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06407_ _02226_ _00074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_241_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07387_ _02612_ soc.spi_video_ram_1.write_fifo.fifo_mem\[29\]\[11\] _03036_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_176_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_182_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09126_ _04294_ _04295_ _00723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_52_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06338_ _02128_ soc.spi_video_ram_1.write_fifo.fifo_mem\[17\]\[4\] _02182_ _02187_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_135_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_191_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_178_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06269_ _02118_ _02141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_09057_ _02116_ _04107_ _02214_ _04257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_108_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_237_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08008_ _02736_ _03646_ _03647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_117_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_219_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_145_wb_clk_i clknet_5_25_0_wb_clk_i clknet_leaf_145_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_46_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_81_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09959_ _04855_ _04848_ _04856_ _00996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_4102 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4113 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4124 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_4135 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_246_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_4146 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4157 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4168 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11921_ _00980_ clknet_leaf_100_wb_clk_i soc.rom_encoder_0.sram_sio_oe vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_185_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_4179 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2700 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_174_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_3445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2711 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2722 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2733 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11852_ _00911_ clknet_leaf_106_wb_clk_i soc.rom_encoder_0.request_data_out\[13\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_57_1400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2744 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2755 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_221_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2766 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10803_ _02231_ soc.spi_video_ram_1.write_fifo.fifo_mem\[7\]\[7\] _05378_ _05386_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_54_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2777 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2788 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_198_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11783_ _00844_ clknet_leaf_104_wb_clk_i soc.rom_encoder_0.output_buffer\[14\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2799 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_207_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_199_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10734_ soc.spi_video_ram_1.write_fifo.fifo_mem\[31\]\[4\] soc.spi_video_ram_1.fifo_in_data\[4\]
+ _05344_ _05349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_10665_ _02219_ soc.spi_video_ram_1.write_fifo.fifo_mem\[29\]\[1\] _05310_ _05312_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_201_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10596_ net17 _05274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_182_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_220_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12335_ _01363_ clknet_leaf_4_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[8\]\[14\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_103_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_182_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_147_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_177_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12266_ _01294_ clknet_leaf_72_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[31\]\[19\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_194_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11217_ _00283_ clknet_leaf_264_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[11\]\[27\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_29_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_123_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput70 net70 io_out[22] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_12197_ _01225_ clknet_leaf_221_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[19\]\[8\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_110_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput81 net81 io_out[8] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_123_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_6060 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11148_ _00214_ clknet_leaf_282_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[14\]\[28\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_110_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6071 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6082 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6093 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_95_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_5370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11079_ _00145_ clknet_leaf_20_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[13\]\[17\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_5381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_231_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_36_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_236_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05640_ _01538_ _01548_ _01549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_64_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3990 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_225_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_1544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_05571_ soc.spi_video_ram_1.output_buffer\[15\] _01475_ _01480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_211_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_205_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_177_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_162_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07310_ _02910_ _02959_ _02960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_176_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08290_ _03837_ _00345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07241_ _02885_ _02887_ _02889_ _02891_ _02892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_34_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_192_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07172_ _02650_ _02825_ _02719_ _02826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_117_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_191_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06123_ _01977_ _01924_ _01990_ _02016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_30_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06054_ _01841_ _01846_ _01947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_191_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_145_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_173_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_207_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_154_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_236_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09813_ soc.rom_encoder_0.request_data_out\[0\] _04743_ _04744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_100_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09744_ _04701_ _00936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_74_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06956_ soc.spi_video_ram_1.write_fifo.fifo_mem\[20\]\[0\] soc.spi_video_ram_1.write_fifo.fifo_mem\[21\]\[0\]
+ soc.spi_video_ram_1.write_fifo.fifo_mem\[22\]\[0\] soc.spi_video_ram_1.write_fifo.fifo_mem\[23\]\[0\]
+ _02591_ _02593_ _02617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_189_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05907_ _01654_ _01802_ _01803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_228_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09675_ _04650_ soc.rom_encoder_0.request_address\[4\] _04632_ _04651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06887_ _02492_ _02551_ _02552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_36_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2007 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2018 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2029 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08626_ _02153_ soc.spi_video_ram_1.write_fifo.fifo_mem\[30\]\[16\] _04011_ _04018_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_199_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05838_ _01595_ _01736_ _01737_ soc.cpu.PC.in\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_203_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08557_ _03981_ _00468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_70_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05769_ _01557_ _01671_ _01672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_168_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07508_ soc.spi_video_ram_1.write_fifo.fifo_mem\[24\]\[26\] soc.spi_video_ram_1.write_fifo.fifo_mem\[25\]\[26\]
+ soc.spi_video_ram_1.write_fifo.fifo_mem\[26\]\[26\] soc.spi_video_ram_1.write_fifo.fifo_mem\[27\]\[26\]
+ _02907_ _02908_ _03156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_146_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_204_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_195_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08488_ _03944_ _00436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_93_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07439_ _02784_ soc.spi_video_ram_1.write_fifo.fifo_mem\[18\]\[27\] _03088_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_11_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10450_ soc.cpu.PC.in\[1\] _05172_ _05173_ _05176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_178_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xcaravel_hack_soc_203 wbs_dat_o[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xcaravel_hack_soc_214 wbs_dat_o[22] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_221_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09109_ _02169_ soc.spi_video_ram_1.write_fifo.fifo_mem\[20\]\[24\] _04258_ _04285_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xcaravel_hack_soc_225 io_oeb[30] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
X_10381_ _02231_ soc.spi_video_ram_1.write_fifo.fifo_mem\[6\]\[7\] _05124_ _05132_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_12120_ _01148_ clknet_leaf_309_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[6\]\[12\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_123_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_12051_ net28 clknet_5_31_0_wb_clk_i soc.rom_encoder_0.data_out\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_215_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_191_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11002_ _00068_ clknet_leaf_265_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[17\]\[27\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_105_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_24_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_218_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11904_ _00963_ clknet_leaf_124_wb_clk_i soc.cpu.DMuxJMP.sel\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_leaf_42_wb_clk_i clknet_5_3_0_wb_clk_i clknet_leaf_42_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_73_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_234_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11835_ _00894_ clknet_leaf_122_wb_clk_i soc.rom_encoder_0.input_buffer\[9\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1840 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1851 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1862 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_158_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1873 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1884 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11766_ _00827_ clknet_leaf_69_wb_clk_i net69 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_144_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1895 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_226_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10717_ _03249_ _05324_ _05339_ _01271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_174_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11697_ _00758_ clknet_leaf_300_wb_clk_i soc.spi_video_ram_1.fifo_in_data\[15\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_9_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_146_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10648_ _05302_ _01239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_173_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10579_ net78 _05261_ _05201_ _05263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_177_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12318_ _01346_ clknet_leaf_115_wb_clk_i soc.ram_encoder_0.data_out\[13\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_115_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12249_ _01277_ clknet_leaf_261_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[31\]\[2\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_155_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_228_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06810_ _02481_ _02485_ _02486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_151_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07790_ _02651_ _03434_ _03435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06741_ _02426_ _00208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_168_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_149_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09460_ soc.rom_encoder_0.output_buffer\[13\] _04504_ _04506_ _02461_ _04507_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_77_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06672_ _02171_ soc.spi_video_ram_1.write_fifo.fifo_mem\[12\]\[25\] _02356_ _02384_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_184_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08411_ soc.spi_video_ram_1.write_fifo.fifo_mem\[27\]\[3\] _02397_ _03899_ _03903_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_240_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05623_ _01467_ soc.spi_video_ram_1.output_buffer\[18\] _01532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_09391_ _01387_ _04453_ soc.spi_video_ram_1.sram_sck_fall_edge _01419_ _04454_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_75_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_178_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08342_ _03865_ _03866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_05554_ soc.spi_video_ram_1.buffer_index\[3\] _01463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_177_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_205_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08273_ soc.ram_encoder_0.output_buffer\[15\] _03814_ _03788_ soc.ram_encoder_0.request_data_out\[11\]
+ _03817_ _03827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_05485_ soc.spi_video_ram_1.write_fifo.write_pointer\[1\] _01400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_193_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_165_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07224_ _02589_ _02875_ _02876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_20_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07155_ _02803_ _02805_ _02807_ _02809_ _02656_ _02810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_195_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06106_ _01902_ _01986_ _01924_ _01998_ _01999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_175_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07086_ _02697_ soc.spi_video_ram_1.write_fifo.fifo_mem\[5\]\[3\] _02742_ _02743_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_105_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_160_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06037_ soc.video_generator_1.v_count\[4\] _01930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_82_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_216_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07988_ soc.spi_video_ram_1.write_fifo.fifo_mem\[20\]\[18\] soc.spi_video_ram_1.write_fifo.fifo_mem\[21\]\[18\]
+ soc.spi_video_ram_1.write_fifo.fifo_mem\[22\]\[18\] soc.spi_video_ram_1.write_fifo.fifo_mem\[23\]\[18\]
+ _02726_ _03041_ _03628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_210_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09727_ _04677_ _04689_ _04690_ _01381_ _00930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_170_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_234_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06939_ _00003_ _02600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_41_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09658_ soc.rom_encoder_0.write_enable _04638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_167_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_216_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08609_ _02136_ soc.spi_video_ram_1.write_fifo.fifo_mem\[30\]\[8\] _04000_ _04009_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_167_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09589_ soc.rom_encoder_0.input_buffer\[4\] _04594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_230_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_169_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_208_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_1414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11620_ _00686_ clknet_leaf_44_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[21\]\[27\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_223_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_169_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11551_ _00617_ clknet_leaf_18_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[25\]\[16\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_184_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_137_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10502_ soc.cpu.PC.REG.data\[11\] soc.cpu.PC.REG.data\[12\] soc.cpu.PC.REG.data\[13\]
+ _05206_ _05215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_32_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11482_ _00548_ clknet_leaf_179_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[24\]\[5\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_leaf_160_wb_clk_i clknet_5_27_0_wb_clk_i clknet_leaf_160_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_155_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10433_ _01589_ _01613_ _01632_ _01652_ _05160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_109_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_164_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10364_ _02114_ _04392_ _05122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_3_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_12103_ _01131_ net85 soc.cpu.ALU.x\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_174_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10295_ _05071_ _05079_ _05080_ _01107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_12034_ _01093_ clknet_leaf_270_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[5\]\[22\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_132_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_232_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_185_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_20_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3050 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3061 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3072 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3083 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_233_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_222_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3094 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11818_ _00877_ clknet_leaf_61_wb_clk_i soc.spi_video_ram_1.write_fifo.read_pointer\[0\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_33_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_248_wb_clk_i clknet_5_19_0_wb_clk_i clknet_leaf_248_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_109_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1692 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11749_ _00810_ clknet_leaf_267_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[4\]\[22\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_175_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_147_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_198_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_198_1749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_200_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_128_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_192_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08960_ _04201_ _00651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_83_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07911_ soc.spi_video_ram_1.write_fifo.fifo_mem\[23\]\[21\] _03554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_130_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08891_ _04164_ _00619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_155_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_229_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07842_ _02607_ _03485_ _03486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_64_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_211_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_216_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07773_ _02924_ soc.spi_video_ram_1.write_fifo.fifo_mem\[6\]\[15\] _03417_ _02895_
+ _03418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_09512_ _02266_ soc.cpu.AReg.data\[8\] _01459_ _04541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06724_ soc.spi_video_ram_1.write_fifo.fifo_mem\[14\]\[14\] _02246_ _02412_ _02418_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_246_1717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09443_ soc.rom_encoder_0.request_data_out\[6\] _03767_ _04493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_06655_ _02375_ _00173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_227_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_212_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_80_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05606_ _01428_ soc.spi_video_ram_1.buffer_index\[5\] _01515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_209_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09374_ soc.spi_video_ram_1.state_sram_clk_counter\[5\] _04441_ _04433_ _04444_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_36_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06586_ soc.spi_video_ram_1.write_fifo.fifo_mem\[13\]\[16\] _02335_ _02328_ _02336_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_33_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08325_ _03855_ _00362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05537_ _01404_ _01446_ _01447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_138_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08256_ _02558_ _03812_ _03813_ _00335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_20_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05468_ soc.spi_video_ram_1.state_counter\[1\] soc.spi_video_ram_1.state_counter\[0\]
+ soc.spi_video_ram_1.state_counter\[3\] soc.spi_video_ram_1.state_counter\[2\] _01384_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_166_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_137_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_192_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07207_ _02710_ _02853_ _02859_ _02606_ _02860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_08187_ _03759_ _00320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_116_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07138_ soc.spi_video_ram_1.write_fifo.fifo_mem\[20\]\[4\] soc.spi_video_ram_1.write_fifo.fifo_mem\[21\]\[4\]
+ soc.spi_video_ram_1.write_fifo.fifo_mem\[22\]\[4\] soc.spi_video_ram_1.write_fifo.fifo_mem\[23\]\[4\]
+ _02717_ _02682_ _02794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_161_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07069_ _02651_ soc.spi_video_ram_1.write_fifo.fifo_mem\[29\]\[2\] _02728_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_216_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5903 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10080_ _04787_ _04934_ _01038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_43_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5914 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5925 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5936 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5947 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5958 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5969 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_235_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10982_ _00048_ clknet_leaf_186_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[17\]\[7\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_112_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_215_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_204_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_231_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_188_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11603_ _00669_ clknet_leaf_20_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[21\]\[10\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_15_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_15_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_11534_ _00600_ clknet_leaf_277_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[23\]\[28\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_54_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_184_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11465_ _00531_ clknet_leaf_20_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[15\]\[17\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_125_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10416_ _02266_ soc.spi_video_ram_1.write_fifo.fifo_mem\[6\]\[24\] _05123_ _05150_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_178_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11396_ _00462_ clknet_leaf_247_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[2\]\[6\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_124_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_193_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_125_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10347_ _01713_ _05103_ _05113_ _01127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_152_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_152_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_239_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10278_ soc.rom_encoder_0.toggled_sram_sck _01396_ _01102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_117_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_215_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12017_ _01076_ clknet_leaf_227_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[5\]\[5\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_78_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_66_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_227_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_93_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_93_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06440_ soc.spi_video_ram_1.write_fifo.fifo_mem\[16\]\[15\] _02248_ _02238_ _02249_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_62_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_221_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_210_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_206_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06371_ _02161_ soc.spi_video_ram_1.write_fifo.fifo_mem\[17\]\[20\] _02181_ _02204_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_222_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08110_ soc.video_generator_1.h_count\[2\] _01990_ _03716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_9_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_175_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09090_ _04275_ _00707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_119_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08041_ _02116_ _01441_ _03677_ _03678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_163_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_190_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_89_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09992_ soc.synch_hack_writeM _01579_ _04880_ _04881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_131_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08943_ soc.spi_video_ram_1.write_fifo.fifo_mem\[22\]\[13\] _04050_ _04189_ _04193_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_83_1462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_233_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_213_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_97_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08874_ soc.spi_video_ram_1.write_fifo.fifo_mem\[25\]\[10\] _02411_ _04155_ _04156_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_215_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3808 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07825_ _02640_ _03463_ _03469_ _03470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_3819 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_217_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_244_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07756_ _03384_ _03391_ _03400_ _03401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_56_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06707_ soc.spi_video_ram_1.fifo_in_data\[8\] _02407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_07687_ _03331_ _03332_ _02577_ _03333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_44_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_213_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09426_ _04473_ _04478_ _04480_ _00839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_77_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06638_ _02366_ _00165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_25_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_197_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_240_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_146_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_181_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09357_ soc.spi_video_ram_1.state_sram_clk_counter\[0\] _04431_ _04432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_06569_ _02326_ _00136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_139_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08308_ _02149_ soc.spi_video_ram_1.write_fifo.fifo_mem\[1\]\[14\] _03842_ _03847_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_205_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09288_ _02214_ _04392_ _04393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_193_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08239_ soc.ram_encoder_0.output_buffer\[11\] _02563_ _03801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_140_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_197_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11250_ _00316_ clknet_leaf_285_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[10\]\[21\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_106_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_238_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_179_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10201_ soc.hack_clock_0.counter\[5\] _05024_ _05026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_136_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11181_ _00247_ clknet_leaf_62_wb_clk_i soc.spi_video_ram_1.output_buffer\[9\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_6401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10132_ _04865_ _04947_ _04948_ _04974_ _04975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_6434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5700 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5711 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5722 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5733 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10063_ _02550_ _04920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_7_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_6489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5744 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_125_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5755 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_212_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_209_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5766 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5777 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5788 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5799 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_169_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_186_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10965_ _00031_ clknet_leaf_67_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[18\]\[19\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_71_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_203_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10896_ _05436_ _01353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_31_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_223_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_156_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11517_ _00583_ clknet_leaf_37_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[23\]\[11\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_172_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11448_ _00514_ clknet_leaf_178_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[15\]\[0\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_125_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_236_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11379_ _00445_ clknet_leaf_30_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[28\]\[18\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_158_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_154_1438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05940_ _01654_ _01833_ _01834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XTAP_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_230_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_79_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05871_ _01595_ _01767_ _01768_ soc.cpu.PC.in\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_15_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_187_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07610_ _02688_ _03256_ _03257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_226_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08590_ _03931_ _02114_ _03998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_leaf_263_wb_clk_i clknet_5_7_0_wb_clk_i clknet_leaf_263_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_35_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_81_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07541_ soc.spi_video_ram_1.write_fifo.fifo_mem\[22\]\[13\] soc.spi_video_ram_1.write_fifo.fifo_mem\[23\]\[13\]
+ _02700_ _03188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_228_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07472_ _02597_ soc.spi_video_ram_1.write_fifo.fifo_mem\[28\]\[12\] _03119_ _02943_
+ _03120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_62_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_34_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_179_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09211_ _00011_ _01752_ _04351_ _00752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_06423_ soc.spi_video_ram_1.fifo_in_data\[10\] _02237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_241_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_163_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09142_ soc.spi_video_ram_1.state_counter\[7\] _04304_ _04306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_148_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06354_ _02195_ _00052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_72_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09073_ _04266_ _00699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_30_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06285_ _02151_ soc.spi_video_ram_1.write_fifo.fifo_mem\[18\]\[15\] _02141_ _02152_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_08024_ _02768_ _03661_ _03662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_163_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_146_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_239_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_1595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_176_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09975_ soc.ram_encoder_0.input_buffer\[9\] _04867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_5007 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_5018 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5029 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08926_ soc.spi_video_ram_1.write_fifo.fifo_mem\[22\]\[5\] _02401_ _04178_ _04184_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_83_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_130_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_213_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_170_1284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08857_ soc.spi_video_ram_1.write_fifo.fifo_mem\[25\]\[2\] _02395_ _04144_ _04147_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_3605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07808_ soc.spi_video_ram_1.write_fifo.fifo_mem\[5\]\[23\] _03453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_3638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2904 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08788_ _04108_ _04109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XTAP_3649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2915 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2926 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2937 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07739_ _02693_ _03380_ _03383_ _02707_ _03384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XTAP_2948 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2959 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_164_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10750_ _05357_ _01286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_240_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_246_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09409_ _02542_ _04464_ _04465_ _04466_ _00836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_129_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_187_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_16_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10681_ _02235_ soc.spi_video_ram_1.write_fifo.fifo_mem\[29\]\[9\] _05310_ _05320_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_90_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_220_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_67_wb_clk_i clknet_5_11_0_wb_clk_i clknet_leaf_67_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_217_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11302_ _00368_ clknet_leaf_297_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[1\]\[28\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12282_ _01310_ clknet_leaf_246_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[7\]\[6\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_135_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_194_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_155_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_11233_ _00299_ clknet_leaf_198_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[10\]\[4\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_107_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_218_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_150_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_6220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_155_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11164_ _00230_ clknet_leaf_149_wb_clk_i soc.ram_encoder_0.output_buffer\[3\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_6231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_171_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10115_ soc.ram_encoder_0.request_data_out\[8\] _04929_ _04962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_67_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_216_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11095_ _00161_ clknet_leaf_260_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[12\]\[4\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_6286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_231_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_5563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10046_ soc.ram_encoder_0.request_address\[9\] soc.ram_encoder_0.address\[9\] _04900_
+ _04909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_29_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4840 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_236_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4851 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4862 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_208_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4873 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4884 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4895 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11997_ _01056_ clknet_leaf_161_wb_clk_i soc.ram_encoder_0.current_state\[0\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_95_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_232_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_229_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10948_ _00014_ clknet_leaf_198_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[18\]\[2\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_32_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_162_1718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_231_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10879_ _01819_ _05221_ _05411_ _05426_ _01346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_242_1753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_220_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_157_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06070_ _01953_ _01957_ _01961_ _01962_ _01963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XANTENNA_1 _01551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_160_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_1243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_193_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_140_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_115_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09760_ _02240_ soc.spi_video_ram_1.write_fifo.fifo_mem\[3\]\[11\] _04708_ _04710_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06972_ _01378_ _02632_ _02633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_112_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_239_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08711_ _03464_ _04046_ _04066_ _00537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_79_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05923_ _01682_ _01812_ _01815_ _01817_ _01818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_09691_ soc.cpu.PC.REG.data\[9\] soc.rom_loader.current_address\[9\] _04638_ _04662_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_39_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08642_ _02169_ soc.spi_video_ram_1.write_fifo.fifo_mem\[30\]\[24\] _03999_ _04026_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_05854_ _01552_ _01717_ soc.cpu.AReg.data\[9\] _01592_ _01753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_132_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_227_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_08573_ _03989_ _00476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05785_ _01685_ _01686_ _01687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_70_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_82_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_07524_ _03167_ _03168_ _03171_ _02706_ _03172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_23_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_222_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07455_ _01419_ _03018_ _03103_ _02677_ _03104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_56_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06406_ soc.spi_video_ram_1.write_fifo.fifo_mem\[16\]\[4\] _02225_ _02217_ _02226_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_210_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07386_ _02924_ soc.spi_video_ram_1.write_fifo.fifo_mem\[30\]\[11\] _02827_ _03035_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_206_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09125_ soc.spi_video_ram_1.state_counter\[1\] soc.spi_video_ram_1.state_counter\[0\]
+ _04295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_194_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06337_ _02186_ _00044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_148_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_198_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09056_ _04256_ _00692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06268_ soc.spi_video_ram_1.fifo_in_data\[10\] _02140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_117_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08007_ soc.spi_video_ram_1.write_fifo.fifo_mem\[24\]\[17\] soc.spi_video_ram_1.write_fifo.fifo_mem\[25\]\[17\]
+ soc.spi_video_ram_1.write_fifo.fifo_mem\[26\]\[17\] soc.spi_video_ram_1.write_fifo.fifo_mem\[27\]\[17\]
+ _02701_ _02737_ _03646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_89_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_135_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_190_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06199_ _01515_ _02076_ _02080_ _02085_ _02086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_144_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_235_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_217_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09958_ net4 _04849_ _04601_ _04856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_131_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_185_wb_clk_i clknet_5_28_0_wb_clk_i clknet_leaf_185_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_4103 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4114 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4125 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08909_ _04173_ _00628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_4136 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_218_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xclkbuf_leaf_114_wb_clk_i clknet_5_26_0_wb_clk_i clknet_leaf_114_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_09889_ _04254_ _04801_ _04803_ _00979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_3402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4147 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4158 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11920_ _00979_ clknet_leaf_99_wb_clk_i net62 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_4169 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2701 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2712 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2723 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11851_ _00910_ clknet_leaf_93_wb_clk_i soc.rom_encoder_0.request_data_out\[12\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_2_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2734 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_167_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2745 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2756 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_214_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10802_ _05385_ _01310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2767 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2778 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11782_ _00843_ clknet_5_14_0_wb_clk_i soc.rom_encoder_0.output_buffer\[13\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2789 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_241_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_198_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10733_ _05348_ _01278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_183_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_213_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_202_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_14_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_224_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10664_ _05311_ _01246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_186_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10595_ _05272_ _05268_ _05273_ _01215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_103_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12334_ _01362_ clknet_leaf_7_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[8\]\[13\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_108_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_177_1246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12265_ _01293_ clknet_leaf_73_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[31\]\[18\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_135_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11216_ _00282_ clknet_leaf_280_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[11\]\[26\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_107_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12196_ _01224_ clknet_leaf_194_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[19\]\[7\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xoutput60 net60 io_out[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput71 net71 io_out[23] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_190_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput82 net82 io_out[9] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_6050 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_151_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11147_ _00213_ clknet_leaf_45_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[14\]\[27\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_6061 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6072 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6083 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6094 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_110_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11078_ _00144_ clknet_leaf_20_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[13\]\[16\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_114_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_23_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_237_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10029_ _04879_ _04900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_209_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_4670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_149_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_110_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4692 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_149_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3980 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3991 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05570_ _01467_ soc.spi_video_ram_1.output_buffer\[14\] _01479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_204_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_177_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07240_ _02650_ _02890_ _02719_ _02891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_73_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_158_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07171_ soc.spi_video_ram_1.write_fifo.fifo_mem\[20\]\[6\] soc.spi_video_ram_1.write_fifo.fifo_mem\[21\]\[6\]
+ soc.spi_video_ram_1.write_fifo.fifo_mem\[22\]\[6\] soc.spi_video_ram_1.write_fifo.fifo_mem\[23\]\[6\]
+ _02645_ _02614_ _02825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_160_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_145_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06122_ _02012_ _02013_ _02014_ _01925_ _02015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_118_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_199_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_201_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_145_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06053_ _01927_ _01938_ _01946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_117_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09812_ _04742_ _04743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_141_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_214_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09743_ _02223_ soc.spi_video_ram_1.write_fifo.fifo_mem\[3\]\[3\] _04697_ _04701_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06955_ _02589_ _02615_ _02616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_246_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05906_ _01669_ _01786_ _01798_ _01801_ _01802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XFILLER_55_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_100_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09674_ soc.cpu.PC.REG.data\[4\] soc.rom_loader.current_address\[4\] _04638_ _04650_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_223_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06886_ _02482_ _02550_ _02551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_27_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2008 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08625_ _04017_ _00500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2019 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05837_ _01552_ _01705_ soc.cpu.AReg.data\[8\] _01592_ _01737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XTAP_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08556_ _02145_ soc.spi_video_ram_1.write_fifo.fifo_mem\[2\]\[12\] _03978_ _03981_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05768_ _01670_ soc.cpu.ALU.x\[5\] _01671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_74_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_242_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_223_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07507_ _02707_ _03147_ _03154_ _02910_ _03155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_19_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08487_ _02138_ soc.spi_video_ram_1.write_fifo.fifo_mem\[28\]\[9\] _03934_ _03944_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_05699_ soc.cpu.ALU.zy _01606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_52_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_168_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07438_ _02691_ _03084_ _03085_ _03086_ _02588_ _03087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_211_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_241_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_195_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07369_ _01964_ _03017_ _02916_ _03018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_6_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xcaravel_hack_soc_204 wbs_dat_o[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_09108_ _04284_ _00716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xcaravel_hack_soc_215 wbs_dat_o[23] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_10380_ _05131_ _01142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_104_1487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xcaravel_hack_soc_226 io_oeb[31] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_202_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09039_ _01408_ _04244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_178_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12050_ net27 clknet_5_31_0_wb_clk_i soc.rom_encoder_0.data_out\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_137_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11001_ _00067_ clknet_leaf_288_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[17\]\[26\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_104_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_172_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_232_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_133_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_8_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_115_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_219_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_133_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11903_ _00962_ clknet_leaf_99_wb_clk_i soc.rom_encoder_0.initialized vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_94_1409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_209_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11834_ _00893_ clknet_leaf_123_wb_clk_i soc.rom_encoder_0.input_buffer\[8\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1830 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_183_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1852 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1863 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_199_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11765_ _00826_ clknet_leaf_69_wb_clk_i soc.spi_video_ram_1.state_sram_clk_counter\[8\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_13_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1874 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_82_wb_clk_i clknet_5_10_0_wb_clk_i clknet_leaf_82_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_1885 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1896 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10716_ soc.spi_video_ram_1.fifo_in_address\[9\] _05325_ _05339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_41_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11696_ _00757_ clknet_leaf_300_wb_clk_i soc.spi_video_ram_1.fifo_in_data\[14\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_leaf_11_wb_clk_i clknet_5_3_0_wb_clk_i clknet_leaf_11_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_201_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10647_ soc.spi_video_ram_1.write_fifo.fifo_mem\[19\]\[22\] _04063_ _05277_ _05302_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_220_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10578_ _01589_ _05261_ _05262_ _01209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_6_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12317_ _01345_ clknet_leaf_114_wb_clk_i soc.ram_encoder_0.data_out\[12\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_157_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_142_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_177_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12248_ _01276_ clknet_leaf_222_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[31\]\[1\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_244_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_218_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12179_ _01207_ clknet_leaf_127_wb_clk_i soc.hack_wait_clocks\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_68_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_231_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06740_ soc.spi_video_ram_1.write_fifo.fifo_mem\[14\]\[22\] _02262_ _02390_ _02426_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_5190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_236_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06671_ _02383_ _00181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_184_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_168_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08410_ _03902_ _00400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05622_ _01468_ _01510_ _01530_ _01531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_18_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09390_ _01388_ _04452_ _04453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_197_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_224_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_205_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_209_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08341_ _03864_ _03865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_162_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05553_ _01461_ soc.spi_video_ram_1.buffer_index\[1\] _01462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_71_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_244_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08272_ _02558_ _03825_ _03826_ _00338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_162_1356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05484_ _01398_ _01399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_123_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07223_ soc.spi_video_ram_1.write_fifo.fifo_mem\[16\]\[8\] soc.spi_video_ram_1.write_fifo.fifo_mem\[17\]\[8\]
+ soc.spi_video_ram_1.write_fifo.fifo_mem\[18\]\[8\] soc.spi_video_ram_1.write_fifo.fifo_mem\[19\]\[8\]
+ _02645_ _02614_ _02875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_164_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_197_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07154_ _02650_ _02808_ _02618_ _02809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_121_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_06105_ _01992_ _01997_ _01923_ _01998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_118_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07085_ _02741_ _02742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_161_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06036_ _01881_ _01855_ _01878_ _01887_ _01929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_47_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_236_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07987_ _02736_ _03626_ _03627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_45_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09726_ net59 _04677_ _04690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06938_ soc.spi_video_ram_1.write_fifo.fifo_mem\[4\]\[0\] soc.spi_video_ram_1.write_fifo.fifo_mem\[5\]\[0\]
+ soc.spi_video_ram_1.write_fifo.fifo_mem\[6\]\[0\] soc.spi_video_ram_1.write_fifo.fifo_mem\[7\]\[0\]
+ _02597_ _02598_ _02599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_21_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_228_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_210_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09657_ _04637_ _00913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06869_ _01654_ _02531_ _02538_ _02539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_2
XFILLER_76_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08608_ _04008_ _00492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09588_ _04592_ _04585_ _04593_ _00888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_187_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08539_ _02128_ soc.spi_video_ram_1.write_fifo.fifo_mem\[2\]\[4\] _03967_ _03972_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_184_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_1448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11550_ _00616_ clknet_leaf_313_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[25\]\[15\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_184_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10501_ _05172_ _05213_ _05214_ _01179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_156_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_7_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11481_ _00547_ clknet_leaf_141_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[24\]\[4\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_183_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_149_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10432_ _01615_ _01802_ _05159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_13_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_221_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10363_ _02539_ _05104_ _05121_ _01135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_48_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_1500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12102_ _01130_ net85 soc.cpu.ALU.x\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_2_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10294_ soc.rom_loader.current_address\[4\] _05078_ _05080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_215_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12033_ _01092_ clknet_leaf_292_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[5\]\[21\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_105_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_24_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_218_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_1353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3040 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3051 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xcaravel_hack_soc_91 io_oeb[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_46_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_3062 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3073 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3084 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_234_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_179_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3095 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_206_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11817_ _00876_ clknet_leaf_60_wb_clk_i soc.spi_video_ram_1.write_fifo.write_pointer\[4\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_128_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_163_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_226_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1693 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11748_ _00809_ clknet_leaf_289_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[4\]\[21\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_230_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_179_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11679_ _00740_ clknet_leaf_63_wb_clk_i soc.video_generator_1.v_count\[7\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_2
Xclkbuf_leaf_288_wb_clk_i clknet_5_4_0_wb_clk_i clknet_leaf_288_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_179_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_239_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_217_wb_clk_i clknet_5_21_0_wb_clk_i clknet_leaf_217_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_115_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_239_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07910_ _02693_ _03549_ _03552_ _02984_ _03553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_237_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08890_ soc.spi_video_ram_1.write_fifo.fifo_mem\[25\]\[18\] _02339_ _04155_ _04164_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_25_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07841_ soc.spi_video_ram_1.write_fifo.fifo_mem\[21\]\[22\] _03485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_190_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_238_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07772_ _02907_ _03416_ _03417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_37_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09511_ _04540_ _00864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06723_ _02417_ _00199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_168_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_237_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_211_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09442_ _04473_ _04491_ _04492_ _00843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_1733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06654_ _02153_ soc.spi_video_ram_1.write_fifo.fifo_mem\[12\]\[16\] _02368_ _02375_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_240_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05605_ _01500_ _01513_ _01514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09373_ soc.spi_video_ram_1.state_sram_clk_counter\[5\] _04441_ _04443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_06585_ soc.spi_video_ram_1.fifo_in_address\[0\] _02335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_205_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08324_ _02165_ soc.spi_video_ram_1.write_fifo.fifo_mem\[1\]\[22\] _03830_ _03855_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_05536_ soc.spi_video_ram_1.write_fifo.write_pointer\[2\] _01445_ _01446_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_178_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_162_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_193_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_1749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08255_ soc.ram_encoder_0.output_buffer\[15\] _02555_ _03813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_220_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_165_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05467_ soc.spi_video_ram_1.state_counter\[5\] soc.spi_video_ram_1.state_counter\[4\]
+ soc.spi_video_ram_1.state_counter\[7\] soc.spi_video_ram_1.state_counter\[6\] _01383_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
X_07206_ _02620_ _02858_ _02859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_105_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08186_ _02171_ soc.spi_video_ram_1.write_fifo.fifo_mem\[10\]\[25\] _03731_ _03759_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_88_1522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07137_ _02678_ _02792_ _02793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_118_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07068_ _02726_ soc.spi_video_ram_1.write_fifo.fifo_mem\[30\]\[2\] _02691_ _02727_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_134_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_161_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06019_ _01836_ _01911_ _01843_ _01912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_88_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5904 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_138_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5915 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5926 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_5937 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5948 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_216_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5959 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_1430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_25_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_229_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09709_ _04674_ soc.rom_encoder_0.request_address\[14\] _04617_ _04675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_10981_ _00047_ clknet_leaf_211_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[17\]\[6\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_5_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_245_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_216_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_1559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_230_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_145_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11602_ _00668_ clknet_leaf_254_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[21\]\[9\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_212_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11533_ _00599_ clknet_leaf_272_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[23\]\[27\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_32_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_144_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11464_ _00530_ clknet_leaf_20_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[15\]\[16\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_172_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_184_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_leaf_310_wb_clk_i clknet_5_0_0_wb_clk_i clknet_leaf_310_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_171_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10415_ _05149_ _01159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_158_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11395_ _00461_ clknet_leaf_212_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[2\]\[5\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_67_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10346_ soc.cpu.ALU.x\[7\] _05109_ _05113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_151_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_140_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_135_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10277_ _04243_ _05067_ _01119_ _01101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_140_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12016_ _01075_ clknet_leaf_254_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[5\]\[4\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_79_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_219_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_150_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_4_0_0_wb_clk_i clknet_3_0_0_wb_clk_i clknet_4_0_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_24_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_222_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_235_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_22_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2180 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06370_ _02203_ _00060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_206_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_202_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_147_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_198_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08040_ _02115_ _01403_ _03677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_200_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_163_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_116_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_192_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_235_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09991_ _04879_ _04880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_143_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08942_ _04192_ _00642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_213_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_229_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_131_1406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08873_ _04142_ _04155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_96_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_245_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07824_ _02952_ _03466_ _03468_ _03469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_3809 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07755_ _02767_ _03392_ _03399_ _02970_ _03400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_37_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06706_ _02406_ _00193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_231_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07686_ _02695_ soc.spi_video_ram_1.write_fifo.fifo_mem\[16\]\[24\] _03332_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_53_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_241_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_198_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_212_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_246_1559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_1563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09425_ soc.rom_encoder_0.output_buffer\[9\] _04479_ _04480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_25_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06637_ _02136_ soc.spi_video_ram_1.write_fifo.fifo_mem\[12\]\[8\] _02357_ _02366_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_129_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06568_ soc.spi_video_ram_1.write_fifo.fifo_mem\[13\]\[8\] _02233_ _02317_ _02326_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_09356_ net69 _04430_ _04431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_200_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_139_wb_clk_i clknet_5_24_0_wb_clk_i clknet_leaf_139_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_127_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08307_ _03846_ _00353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_90_1478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05519_ soc.spi_video_ram_1.state_sram_clk_counter\[7\] _01432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_09287_ soc.spi_video_ram_1.write_fifo.write_pointer\[4\] _01403_ _03862_ _04392_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_139_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06499_ _02134_ soc.spi_video_ram_1.write_fifo.fifo_mem\[0\]\[7\] _02279_ _02287_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_107_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08238_ soc.ram_encoder_0.output_buffer\[7\] _03781_ _03789_ soc.ram_encoder_0.request_data_out\[3\]
+ _03799_ _03800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_176_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_222_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08169_ _03750_ _00311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_134_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10200_ _05017_ _05024_ _05025_ _01068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_180_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11180_ _00246_ clknet_leaf_58_wb_clk_i soc.spi_video_ram_1.output_buffer\[10\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_133_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10131_ soc.ram_encoder_0.request_data_out\[12\] _04929_ _04974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_6424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_122_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5701 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_47_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_1514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_6446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_7_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_6457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5712 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_88_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5723 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10062_ _02112_ _02499_ _04919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_6479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5734 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_173_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5745 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_197_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5756 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5767 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_87_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5778 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5789 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_235_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_188_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_204_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_217_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10964_ _00030_ clknet_leaf_76_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[18\]\[18\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_182_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_231_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_188_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10895_ soc.spi_video_ram_1.write_fifo.fifo_mem\[8\]\[4\] soc.spi_video_ram_1.fifo_in_data\[4\]
+ _05431_ _05436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_70_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_240_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_145_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11516_ _00582_ clknet_leaf_14_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[23\]\[10\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_201_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_141_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12496_ net57 net56 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_8_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11447_ _00513_ clknet_leaf_302_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[30\]\[28\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_153_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_193_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11378_ _00444_ clknet_leaf_73_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[28\]\[17\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_4_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_217_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10329_ _05102_ _05103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_227_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05870_ _01552_ _01702_ soc.cpu.AReg.data\[10\] _01591_ _01768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_187_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07540_ _03015_ _03186_ _03187_ _00245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_223_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07471_ _02931_ _03118_ _03119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_165_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_210_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06422_ _02236_ _00079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09210_ soc.spi_video_ram_1.fifo_in_data\[9\] _04346_ _04351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_206_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_232_wb_clk_i clknet_5_5_0_wb_clk_i clknet_leaf_232_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_09141_ _04294_ _04304_ _04305_ _00728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_33_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06353_ _02143_ soc.spi_video_ram_1.write_fifo.fifo_mem\[17\]\[11\] _02193_ _02195_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_09072_ _02229_ soc.spi_video_ram_1.write_fifo.fifo_mem\[20\]\[6\] _04259_ _04266_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06284_ soc.spi_video_ram_1.fifo_in_data\[15\] _02151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_135_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08023_ soc.spi_video_ram_1.write_fifo.fifo_mem\[8\]\[16\] soc.spi_video_ram_1.write_fifo.fifo_mem\[9\]\[16\]
+ soc.spi_video_ram_1.write_fifo.fifo_mem\[10\]\[16\] soc.spi_video_ram_1.write_fifo.fifo_mem\[11\]\[16\]
+ _02769_ _02770_ _03661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_129_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_190_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_162_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_116_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_172_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_171_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09974_ _04865_ _04848_ _04866_ _01001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_5008 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5019 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08925_ _04183_ _00634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_170_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_4318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08856_ _04146_ _00602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_131_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_217_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07807_ _02920_ soc.spi_video_ram_1.write_fifo.fifo_mem\[6\]\[23\] _03451_ _02838_
+ _03452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_3628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05999_ soc.video_generator_1.h_count\[3\] soc.video_generator_1.h_count\[4\] _01842_
+ _01892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08787_ _02116_ _01445_ _04107_ _04108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_2905 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2916 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2927 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07738_ _03381_ _03382_ _02976_ _03383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_2938 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_169_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2949 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_213_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_246_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_183_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_38_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_246_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07669_ _02573_ soc.spi_video_ram_1.write_fifo.fifo_mem\[12\]\[14\] _03315_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_129_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_186_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_197_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09408_ soc.rom_encoder_0.request_address\[5\] _02543_ _04466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_129_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_186_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10680_ _05319_ _01254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_55_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_201_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_179_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09339_ _04420_ _00811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_107_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_205_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_187_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_193_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_194_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11301_ _00367_ clknet_leaf_43_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[1\]\[27\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12281_ _01309_ clknet_leaf_245_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[7\]\[5\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_112_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_14_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_181_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11232_ _00298_ clknet_leaf_260_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[10\]\[3\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_84_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_150_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11163_ _00229_ clknet_leaf_149_wb_clk_i soc.ram_encoder_0.output_buffer\[4\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_6210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_36_wb_clk_i clknet_5_2_0_wb_clk_i clknet_leaf_36_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_6232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_122_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_6243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10114_ _04952_ _04961_ _01045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_6254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_136_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11094_ _00160_ clknet_leaf_261_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[12\]\[3\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_6265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_212_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_209_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_118_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10045_ _04908_ _01030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_27_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4830 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4841 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4852 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_4863 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4874 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4885 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_4896 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_205_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11996_ _01055_ clknet_leaf_161_wb_clk_i soc.ram_encoder_0.sram_sio_oe vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_17_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_21_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_189_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_186_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10947_ _00013_ clknet_leaf_216_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[18\]\[1\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_44_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10878_ soc.ram_encoder_0.data_out\[13\] _05426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_223_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_203_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_185_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_157_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_172_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_145_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_2 _02856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_160_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_236_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_141_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_154_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_1591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06971_ soc.spi_video_ram_1.current_state\[0\] _01411_ _02629_ _02630_ _02631_ _02632_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_4
XFILLER_230_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_171_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08710_ _04065_ _04048_ _04066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_05922_ _01682_ _01816_ _01817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09690_ _04661_ _00922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_80_1477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05853_ _01654_ _01751_ _01752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_08641_ _04025_ _00508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_81_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_242_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_187_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05784_ _01598_ soc.cpu.AReg.data\[6\] _01606_ _01686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_08572_ _02161_ soc.spi_video_ram_1.write_fifo.fifo_mem\[2\]\[20\] _03966_ _03989_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XPHY_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_54_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_228_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_169_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07523_ _02763_ soc.spi_video_ram_1.write_fifo.fifo_mem\[14\]\[26\] _03170_ _02592_
+ _03171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_63_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_211_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_179_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_168_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07454_ _03063_ _03102_ _03103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06405_ soc.spi_video_ram_1.fifo_in_data\[4\] _02225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_50_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07385_ _02696_ soc.spi_video_ram_1.write_fifo.fifo_mem\[31\]\[11\] _03034_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_148_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06336_ _02126_ soc.spi_video_ram_1.write_fifo.fifo_mem\[17\]\[3\] _02182_ _02186_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_09124_ soc.spi_video_ram_1.state_counter\[0\] _04294_ _00722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_202_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_175_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09055_ _04254_ _04255_ _04256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_06267_ _02139_ _00021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_191_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08006_ _03638_ _03640_ _03642_ _03644_ _02710_ _03645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_191_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06198_ _02074_ _02082_ _02083_ _02084_ _02085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_117_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09957_ soc.ram_encoder_0.input_buffer\[3\] _04855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_4104 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_213_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4115 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08908_ soc.spi_video_ram_1.write_fifo.fifo_mem\[25\]\[27\] _02351_ _04143_ _04173_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_115_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09888_ _04738_ _04800_ _04802_ _04803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XTAP_4126 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4137 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4148 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4159 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08839_ _03431_ _04124_ _04136_ _00595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_98_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_246_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_245_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2702 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2713 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11850_ _00909_ clknet_leaf_107_wb_clk_i soc.rom_encoder_0.request_data_out\[11\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_22_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2724 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2735 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_154_wb_clk_i clknet_5_30_0_wb_clk_i clknet_leaf_154_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_2746 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10801_ _02229_ soc.spi_video_ram_1.write_fifo.fifo_mem\[7\]\[6\] _05378_ _05385_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_2757 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_26_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2768 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11781_ _00842_ clknet_leaf_104_wb_clk_i soc.rom_encoder_0.output_buffer\[12\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2779 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_226_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_144_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_148_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10732_ soc.spi_video_ram_1.write_fifo.fifo_mem\[31\]\[3\] soc.spi_video_ram_1.fifo_in_data\[3\]
+ _05344_ _05348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_242_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10663_ _02213_ soc.spi_video_ram_1.write_fifo.fifo_mem\[29\]\[0\] _05310_ _05311_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_139_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_220_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_167_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_167_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10594_ soc.gpio_i_stored\[2\] _05268_ _02053_ _05273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_51_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_12333_ _01361_ clknet_leaf_2_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[8\]\[12\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_33_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12264_ _01292_ clknet_leaf_73_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[31\]\[17\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_123_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_218_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11215_ _00281_ clknet_leaf_236_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[11\]\[25\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12195_ _01223_ clknet_leaf_247_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[19\]\[6\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xoutput50 net50 io_oeb[16] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput61 net61 io_out[13] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_150_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput72 net72 io_out[24] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_6040 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11146_ _00212_ clknet_leaf_278_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[14\]\[26\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xoutput83 net83 la_data_out[27] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_6051 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6062 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_231_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6073 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6084 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_7_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11077_ _00143_ clknet_leaf_3_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[13\]\[15\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_6095 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_236_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10028_ _04899_ _01022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_114_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_23_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4693 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_224_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3970 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_52_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3981 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_1513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_229_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3992 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11979_ _01038_ clknet_leaf_157_wb_clk_i soc.ram_data_out\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_17_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_166_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_220_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07170_ _02589_ _02823_ _02824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_157_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_203_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06121_ _01976_ _01991_ _02014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_173_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06052_ _01927_ _01938_ _01944_ _01945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_133_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_193_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09811_ _04567_ _04742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_140_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_115_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_246_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_228_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09742_ _04700_ _00935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_41_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06954_ soc.spi_video_ram_1.write_fifo.fifo_mem\[16\]\[0\] soc.spi_video_ram_1.write_fifo.fifo_mem\[17\]\[0\]
+ soc.spi_video_ram_1.write_fifo.fifo_mem\[18\]\[0\] soc.spi_video_ram_1.write_fifo.fifo_mem\[19\]\[0\]
+ _02613_ _02614_ _02615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_101_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_210_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05905_ _01799_ _01800_ _01796_ _01669_ _01801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_09673_ _04618_ _04648_ _04649_ _00917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06885_ soc.ram_encoder_0.initializing_step\[2\] soc.ram_encoder_0.initializing_step\[1\]
+ _02549_ _02550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_132_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_227_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2009 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08624_ _02151_ soc.spi_video_ram_1.write_fifo.fifo_mem\[30\]\[15\] _04011_ _04017_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_94_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05836_ _01654_ _01735_ _01736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_243_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_184_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08555_ _03980_ _00467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05767_ _01558_ _01670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_145_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_93_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07506_ _02588_ _03150_ _03153_ _03154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_126_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_208_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_165_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05698_ _01601_ _01573_ _01602_ _01604_ _01579_ _01605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_08486_ _03943_ _00435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_243_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_196_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07437_ _02922_ soc.spi_video_ram_1.write_fifo.fifo_mem\[23\]\[27\] _02722_ _03086_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_210_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_4_13_0_wb_clk_i clknet_3_6_0_wb_clk_i clknet_4_13_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_149_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_206_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_221_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07368_ _01939_ _02034_ _03017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_143_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09107_ _02167_ soc.spi_video_ram_1.write_fifo.fifo_mem\[20\]\[23\] _04258_ _04284_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_52_1398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xcaravel_hack_soc_205 wbs_dat_o[13] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_164_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06319_ _02174_ _00038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_164_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xcaravel_hack_soc_216 wbs_dat_o[24] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_07299_ _02597_ soc.spi_video_ram_1.write_fifo.fifo_mem\[17\]\[10\] _02949_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xcaravel_hack_soc_227 io_oeb[32] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_108_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_184_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09038_ _01378_ _04243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_190_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_219_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11000_ _00066_ clknet_leaf_235_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[17\]\[25\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_104_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_131_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_218_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_150_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11902_ _00961_ clknet_leaf_296_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[3\]\[28\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_206_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11833_ _00892_ clknet_leaf_122_wb_clk_i soc.rom_encoder_0.input_buffer\[7\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_27_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_233_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1820 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1831 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1842 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_198_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1853 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_183_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1864 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11764_ _00825_ clknet_leaf_68_wb_clk_i soc.spi_video_ram_1.state_sram_clk_counter\[7\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffnq_2
XTAP_1875 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_202_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1886 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10715_ _03347_ _05324_ _05338_ _01270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_1897 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11695_ _00756_ clknet_leaf_301_wb_clk_i soc.spi_video_ram_1.fifo_in_data\[13\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_186_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10646_ _05301_ _01238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_70_1465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_167_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_155_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10577_ net77 _05261_ _05201_ _05262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xclkbuf_leaf_51_wb_clk_i clknet_5_6_0_wb_clk_i clknet_leaf_51_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_122_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_196_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12316_ _01344_ clknet_leaf_117_wb_clk_i soc.ram_encoder_0.data_out\[11\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_127_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12247_ _01275_ clknet_leaf_187_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[31\]\[0\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_68_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_190_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_12178_ _01206_ clknet_5_15_0_wb_clk_i soc.rom_encoder_0.write_enable vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_151_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_151_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11129_ _00195_ clknet_leaf_201_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[14\]\[9\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_27_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_237_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5180 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_209_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06670_ _02169_ soc.spi_video_ram_1.write_fifo.fifo_mem\[12\]\[24\] _02356_ _02383_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_64_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_149_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_225_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_188_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_184_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_97_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_184_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_05621_ _01467_ soc.spi_video_ram_1.output_buffer\[17\] _01530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_64_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_184_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_149_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08340_ _02388_ _03863_ _03864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05552_ soc.spi_video_ram_1.buffer_index\[0\] _01461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_127_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08271_ soc.ram_encoder_0.output_buffer\[18\] _02555_ _03826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_33_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_225_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05483_ soc.spi_video_ram_1.write_fifo.read_pointer\[2\] soc.spi_video_ram_1.write_fifo.write_pointer\[2\]
+ _01398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_127_1477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_20_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_207_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07222_ _02583_ _02873_ _02640_ _02874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_34_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_146_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07153_ soc.spi_video_ram_1.write_fifo.fifo_mem\[4\]\[5\] soc.spi_video_ram_1.write_fifo.fifo_mem\[5\]\[5\]
+ soc.spi_video_ram_1.write_fifo.fifo_mem\[6\]\[5\] soc.spi_video_ram_1.write_fifo.fifo_mem\[7\]\[5\]
+ _02651_ _02652_ _02808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_118_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_199_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06104_ _01989_ _01993_ _01996_ _01925_ _01997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_161_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07084_ _02740_ _02741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_173_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_172_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06035_ _01881_ _01855_ _01928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_133_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_214_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07986_ soc.spi_video_ram_1.write_fifo.fifo_mem\[16\]\[18\] soc.spi_video_ram_1.write_fifo.fifo_mem\[17\]\[18\]
+ soc.spi_video_ram_1.write_fifo.fifo_mem\[18\]\[18\] soc.spi_video_ram_1.write_fifo.fifo_mem\[19\]\[18\]
+ _02701_ _03041_ _03626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_25_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09725_ soc.ram_encoder_0.output_buffer\[17\] _03814_ _03788_ soc.ram_encoder_0.request_data_out\[13\]
+ _03817_ _04689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_170_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_74_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06937_ _02592_ _02598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_60_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09656_ soc.rom_encoder_0.data_out\[15\] soc.rom_encoder_0.request_data_out\[15\]
+ _04632_ _04637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_41_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_167_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06868_ _02534_ _02536_ _02537_ _02538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_28_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08607_ _02134_ soc.spi_video_ram_1.write_fifo.fifo_mem\[30\]\[7\] _04000_ _04008_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_215_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05819_ _01618_ soc.cpu.AReg.data\[8\] _01718_ soc.ram_data_out\[8\] _01719_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_09587_ net8 _04586_ _04553_ _04593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06799_ net67 _02453_ _02476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_242_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08538_ _03971_ _00459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_58_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_180_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08469_ _02113_ soc.spi_video_ram_1.write_fifo.fifo_mem\[28\]\[0\] _03934_ _03935_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_211_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10500_ soc.cpu.PC.in\[13\] _05188_ _05201_ _05214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_17_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11480_ _00546_ clknet_leaf_141_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[24\]\[3\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_195_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10431_ _01615_ _01766_ _05158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
Xclkbuf_5_2_0_wb_clk_i clknet_4_1_0_wb_clk_i clknet_5_2_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_109_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_192_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10362_ soc.cpu.ALU.x\[15\] _05102_ _05121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_139_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_178_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_174_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_191_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12101_ _01129_ net85 soc.cpu.ALU.x\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10293_ soc.rom_loader.current_address\[4\] _05078_ _05079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_139_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12032_ _01091_ clknet_leaf_59_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[5\]\[20\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_104_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_191_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_219_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_93_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_3030 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_207_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3041 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3052 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_189_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xcaravel_hack_soc_92 io_oeb[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_3063 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3074 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3085 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3096 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11816_ _00875_ clknet_leaf_48_wb_clk_i soc.spi_video_ram_1.write_fifo.write_pointer\[3\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_18_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_199_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1694 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11747_ _00808_ clknet_leaf_59_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[4\]\[20\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_14_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_187_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_187_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11678_ _00739_ clknet_leaf_64_wb_clk_i soc.video_generator_1.v_count\[6\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_204_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_190_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10629_ soc.spi_video_ram_1.write_fifo.fifo_mem\[19\]\[13\] _04050_ _05289_ _05293_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_128_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_183_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_170_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_154_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_170_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_170_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_257_wb_clk_i clknet_5_18_0_wb_clk_i clknet_leaf_257_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_64_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_97_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07840_ _02764_ soc.spi_video_ram_1.write_fifo.fifo_mem\[22\]\[22\] _03483_ _02958_
+ _03484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_57_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_231_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07771_ soc.spi_video_ram_1.write_fifo.fifo_mem\[7\]\[15\] _03416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_42_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09510_ _02264_ soc.cpu.AReg.data\[7\] _04339_ _04540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_83_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06722_ soc.spi_video_ram_1.write_fifo.fifo_mem\[14\]\[13\] _02244_ _02412_ _02417_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_1701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09441_ soc.rom_encoder_0.output_buffer\[13\] _04479_ _04492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_37_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06653_ _02374_ _00172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_1745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_55_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_224_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_168_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05604_ soc.spi_video_ram_1.buffer_index\[4\] _01488_ _01506_ _01512_ _01513_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_09372_ _04441_ _04442_ _00822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_36_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06584_ _02334_ _00143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_244_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_240_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08323_ _03854_ _00361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_55_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05535_ _01400_ _01444_ _01445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_127_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_222_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08254_ soc.ram_encoder_0.request_address\[14\] _02506_ _03789_ soc.ram_encoder_0.request_data_out\[7\]
+ _03811_ _03812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_123_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05466_ soc.spi_video_ram_1.state_counter\[9\] soc.spi_video_ram_1.state_counter\[8\]
+ soc.spi_video_ram_1.state_counter\[10\] _01382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_197_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07205_ _02854_ _02855_ _02856_ _02857_ _02570_ _02719_ _02858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_08185_ _03758_ _00319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_119_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_229_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_174_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_146_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07136_ soc.spi_video_ram_1.write_fifo.fifo_mem\[16\]\[4\] soc.spi_video_ram_1.write_fifo.fifo_mem\[17\]\[4\]
+ soc.spi_video_ram_1.write_fifo.fifo_mem\[18\]\[4\] soc.spi_video_ram_1.write_fifo.fifo_mem\[19\]\[4\]
+ _02681_ _02758_ _02792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_146_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07067_ _02607_ _02726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_106_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06018_ _01837_ _01839_ _01911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_5905 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_173_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5916 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5927 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5938 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5949 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07969_ _03577_ _03609_ _03579_ _03610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_21_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_228_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09708_ soc.cpu.PC.REG.data\[14\] soc.rom_loader.current_address\[14\] _04638_ _04674_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_210_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10980_ _00046_ clknet_leaf_226_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[17\]\[5\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_95_1505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_244_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09639_ soc.rom_encoder_0.data_out\[7\] soc.rom_encoder_0.request_data_out\[7\] _04621_
+ _04628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_15_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_147_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_243_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11601_ _00667_ clknet_leaf_207_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[21\]\[8\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_142_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_145_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_230_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_208_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11532_ _00598_ clknet_leaf_281_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[23\]\[26\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_183_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11463_ _00529_ clknet_leaf_9_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[15\]\[15\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_221_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10414_ _02264_ soc.spi_video_ram_1.write_fifo.fifo_mem\[6\]\[23\] _05123_ _05149_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_165_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11394_ _00460_ clknet_leaf_198_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[2\]\[4\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_136_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10345_ _01699_ _05103_ _05112_ _01126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_174_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_155_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_140_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10276_ _05068_ _01119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_105_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_234_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12015_ _01074_ clknet_leaf_265_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[5\]\[3\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_66_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_187_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_165_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_34_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_59_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_234_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_185_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_206_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_245_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2170 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2181 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_222_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_226_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_175_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_156_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_200_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09990_ _04831_ _04878_ _04879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_143_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_131_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08941_ soc.spi_video_ram_1.write_fifo.fifo_mem\[22\]\[12\] _04047_ _04189_ _04192_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_103_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_237_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_174_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08872_ _04154_ _00610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_85_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_131_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07823_ _02704_ soc.spi_video_ram_1.write_fifo.fifo_mem\[13\]\[23\] _03467_ _02742_
+ _03468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_69_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_229_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07754_ _02582_ _03395_ _03398_ _03399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_22_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_226_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_211_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06705_ soc.spi_video_ram_1.write_fifo.fifo_mem\[14\]\[7\] _02405_ _02391_ _02406_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_07685_ _02783_ soc.spi_video_ram_1.write_fifo.fifo_mem\[17\]\[24\] _03331_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_25_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09424_ _02541_ _04479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_225_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06636_ _02365_ _00164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_90_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_205_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_241_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09355_ soc.spi_video_ram_1.state_counter\[0\] _04428_ _04429_ _04430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_100_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06567_ _02325_ _00135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_212_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08306_ _02147_ soc.spi_video_ram_1.write_fifo.fifo_mem\[1\]\[13\] _03842_ _03846_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_51_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05518_ _01429_ _01431_ _01396_ _00008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_139_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09286_ _04391_ _00787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_166_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_165_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06498_ _02286_ _00105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08237_ soc.ram_encoder_0.request_address\[10\] _02505_ _03799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_14_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_179_wb_clk_i clknet_5_23_0_wb_clk_i clknet_leaf_179_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_147_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08168_ _02153_ soc.spi_video_ram_1.write_fifo.fifo_mem\[10\]\[16\] _03743_ _03750_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_118_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_108_wb_clk_i clknet_5_15_0_wb_clk_i clknet_leaf_108_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_134_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07119_ soc.spi_video_ram_1.write_fifo.fifo_mem\[0\]\[4\] soc.spi_video_ram_1.write_fifo.fifo_mem\[1\]\[4\]
+ soc.spi_video_ram_1.write_fifo.fifo_mem\[2\]\[4\] soc.spi_video_ram_1.write_fifo.fifo_mem\[3\]\[4\]
+ _02713_ _02714_ _02775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_101_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08099_ soc.spi_video_ram_1.write_fifo.fifo_mem\[11\]\[27\] _02351_ _03679_ _03709_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_134_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_192_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_171_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10130_ _04952_ _04973_ _01049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_6414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_238_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_106_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_192_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_6447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5702 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5713 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10061_ _04917_ _04918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_5724 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_134_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_216_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5735 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5746 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5757 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5768 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_130_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5779 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_229_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_169_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_229_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10963_ _00029_ clknet_leaf_79_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[18\]\[17\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_216_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_229_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10894_ _05435_ _01352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_204_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_227_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_231_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_145_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_196_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_157_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11515_ _00581_ clknet_leaf_253_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[23\]\[9\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_102_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_200_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12495_ net57 net55 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_172_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_184_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11446_ _00512_ clknet_leaf_41_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[30\]\[27\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_165_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_201_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11377_ _00443_ clknet_leaf_30_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[28\]\[16\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_140_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10328_ _01553_ soc.cpu.instruction\[4\] _05102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XTAP_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10259_ soc.spi_video_ram_1.fifo_in_address\[8\] _05045_ _05058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_67_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_113_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_187_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_208_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_241_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_235_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_207_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07470_ soc.spi_video_ram_1.write_fifo.fifo_mem\[29\]\[12\] _03118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_78_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_223_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_201_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06421_ soc.spi_video_ram_1.write_fifo.fifo_mem\[16\]\[9\] _02235_ _02217_ _02236_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_72_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09140_ soc.spi_video_ram_1.state_counter\[6\] _04302_ _04305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_06352_ _02194_ _00051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_33_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_6_wb_clk_i clknet_5_0_0_wb_clk_i clknet_leaf_6_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_147_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_198_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_206_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06283_ _02150_ _00026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09071_ _04265_ _00698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_124_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_163_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_272_wb_clk_i clknet_5_6_0_wb_clk_i clknet_leaf_272_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_163_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08022_ _03577_ _03659_ _02720_ _03660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_144_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_201_wb_clk_i clknet_5_19_0_wb_clk_i clknet_leaf_201_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_235_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_157_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09973_ soc.ram_encoder_0.input_buffer\[4\] _04847_ _04248_ _04866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_130_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5009 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08924_ soc.spi_video_ram_1.write_fifo.fifo_mem\[22\]\[4\] _02399_ _04178_ _04183_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_135_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_135_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08855_ soc.spi_video_ram_1.write_fifo.fifo_mem\[25\]\[1\] _02393_ _04144_ _04146_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_97_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07806_ _02688_ _03450_ _03451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_84_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08786_ _02115_ _01403_ _04107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_05998_ soc.video_generator_1.h_count\[3\] _01842_ _01891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_26_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_233_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2906 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2917 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07737_ _02922_ soc.spi_video_ram_1.write_fifo.fifo_mem\[16\]\[15\] _03382_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2928 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2939 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_198_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07668_ _02931_ soc.spi_video_ram_1.write_fifo.fifo_mem\[14\]\[14\] _03313_ _02646_
+ _03314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_25_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09407_ soc.rom_encoder_0.output_buffer\[6\] _02541_ _04465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06619_ _02355_ _02356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_07599_ soc.spi_video_ram_1.write_fifo.fifo_mem\[31\]\[25\] _03246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_200_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_213_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09338_ _02264_ soc.spi_video_ram_1.write_fifo.fifo_mem\[4\]\[23\] _04394_ _04420_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_51_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_178_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09269_ _02258_ soc.spi_video_ram_1.write_fifo.fifo_mem\[9\]\[20\] _04359_ _04383_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_103_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11300_ _00366_ clknet_leaf_293_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[1\]\[26\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_166_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_153_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_12280_ _01308_ clknet_leaf_258_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[7\]\[4\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_119_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11231_ _00297_ clknet_leaf_137_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[10\]\[2\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_4_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_150_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_135_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11162_ _00228_ clknet_leaf_92_wb_clk_i soc.rom_encoder_0.output_buffer\[1\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_155_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_6211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_6233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_171_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10113_ soc.ram_data_out\[7\] _04927_ _04960_ _04961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_96_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11093_ _00159_ clknet_leaf_54_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[12\]\[2\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_6266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_49_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_6288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10044_ soc.ram_encoder_0.request_address\[8\] soc.ram_encoder_0.address\[8\] _04900_
+ _04908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_5565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4820 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_76_wb_clk_i clknet_5_8_0_wb_clk_i clknet_leaf_76_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_5576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4831 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_102_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4842 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4853 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4864 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4875 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4886 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4897 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_223_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11995_ _01054_ clknet_leaf_161_wb_clk_i net81 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_16_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_217_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_95_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_182_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10946_ _00012_ clknet_leaf_207_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[18\]\[0\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_32_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_225_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_205_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_1430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10877_ _01803_ _05221_ _05411_ _05425_ _01345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_143_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_31_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_203_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_129_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_125_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_185_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_199_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_3 _02907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11429_ _00495_ clknet_leaf_11_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[30\]\[10\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_154_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_141_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06970_ soc.spi_video_ram_1.current_state\[4\] _01417_ _01391_ _02631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_100_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05921_ _01807_ _01810_ _01816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_20_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08640_ _02167_ soc.spi_video_ram_1.write_fifo.fifo_mem\[30\]\[23\] _03999_ _04025_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_66_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05852_ _01682_ _01748_ _01749_ _01750_ _01751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_55_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_215_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_212_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08571_ _03988_ _00475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05783_ soc.ram_data_out\[6\] _01579_ _01573_ net43 _01563_ _01685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_35_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_07522_ _02590_ _03169_ _03170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_81_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07453_ _02918_ _03082_ _03101_ _03102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_62_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06404_ _02224_ _00073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_195_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07384_ soc.spi_video_ram_1.write_fifo.fifo_mem\[24\]\[11\] soc.spi_video_ram_1.write_fifo.fifo_mem\[25\]\[11\]
+ soc.spi_video_ram_1.write_fifo.fifo_mem\[26\]\[11\] soc.spi_video_ram_1.write_fifo.fifo_mem\[27\]\[11\]
+ _02688_ _02827_ _03033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_37_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09123_ _04293_ _04294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_06335_ _02185_ _00043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_176_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_148_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09054_ soc.spi_video_ram_1.write_fifo.read_pointer\[4\] _04253_ _04255_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_178_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06266_ _02138_ soc.spi_video_ram_1.write_fifo.fifo_mem\[18\]\[9\] _02120_ _02139_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_190_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_159_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_194_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_159_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08005_ _02685_ _03643_ _02720_ _03644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_191_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_237_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06197_ _01517_ _01519_ _02084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_104_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_172_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_89_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09956_ _04853_ _04848_ _04854_ _00995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_63_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08907_ _04172_ _00627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_246_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4105 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_170_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09887_ _02438_ _04730_ _02450_ _02444_ _04802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XTAP_4116 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_4127 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_131_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4138 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4149 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08838_ _04065_ _04110_ _04136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_3404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_230_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_131_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2703 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2714 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_205_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08769_ _04098_ _00563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_113_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2725 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2736 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_199_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10800_ _05384_ _01309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2747 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2758 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_183_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11780_ _00841_ clknet_leaf_104_wb_clk_i soc.rom_encoder_0.output_buffer\[11\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_2769 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10731_ _05347_ _01277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_207_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_186_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_201_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xclkbuf_leaf_194_wb_clk_i clknet_5_25_0_wb_clk_i clknet_leaf_194_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_10662_ _05309_ _05310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_185_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_123_wb_clk_i clknet_5_15_0_wb_clk_i clknet_leaf_123_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_107_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_222_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10593_ net16 _05272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_12332_ _01360_ clknet_leaf_42_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[8\]\[11\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_31_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_177_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_181_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12263_ _01291_ clknet_leaf_26_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[31\]\[16\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_107_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11214_ _00280_ clknet_leaf_304_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[11\]\[24\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_123_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12194_ _01222_ clknet_leaf_217_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[19\]\[5\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_123_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput51 net51 io_oeb[17] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_155_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput62 net62 io_out[14] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_6030 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput73 net73 io_out[25] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_11145_ _00211_ clknet_leaf_285_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[14\]\[25\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_6041 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_110_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6052 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6063 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6074 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6085 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11076_ _00142_ clknet_leaf_5_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[13\]\[14\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_6096 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_49_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10027_ soc.ram_encoder_0.request_address\[0\] soc.ram_encoder_0.address\[0\] _04889_
+ _04899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_3_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_4683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_149_1317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_4694 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3960 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3971 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3982 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3993 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_189_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11978_ _01037_ clknet_leaf_127_wb_clk_i soc.ram_encoder_0.initialized vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_63_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10929_ _05453_ _01369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_147_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_158_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_158_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_242_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06120_ _01986_ _01924_ _01991_ _02013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_9_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_117_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_173_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_172_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_195_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06051_ _01942_ _01943_ _01944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_114_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_236_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_160_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09810_ _04739_ _04741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_98_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09741_ _02221_ soc.spi_video_ram_1.write_fifo.fifo_mem\[3\]\[2\] _04697_ _04700_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_154_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06953_ _02592_ _02614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_3
X_05904_ _01793_ _01794_ _01800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_09672_ soc.rom_encoder_0.request_address\[3\] _04618_ _04649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_55_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06884_ soc.ram_encoder_0.initializing_step\[4\] soc.ram_encoder_0.initializing_step\[3\]
+ _02549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_132_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_228_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08623_ _04016_ _00499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_05835_ _01669_ _01722_ _01731_ _01734_ _01735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_3_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_242_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08554_ _02143_ soc.spi_video_ram_1.write_fifo.fifo_mem\[2\]\[11\] _03978_ _03980_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_05766_ _01585_ _01669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_51_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07505_ _02744_ soc.spi_video_ram_1.write_fifo.fifo_mem\[22\]\[26\] _03152_ _02908_
+ _03153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_39_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_211_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_168_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08485_ _02136_ soc.spi_video_ram_1.write_fifo.fifo_mem\[28\]\[8\] _03934_ _03943_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_05697_ soc.gpio_i_stored\[1\] _01564_ _01603_ _01576_ _01604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_51_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_39_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07436_ _02752_ soc.spi_video_ram_1.write_fifo.fifo_mem\[22\]\[27\] _03085_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_50_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_167_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07367_ _03014_ _03015_ _03016_ _00243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_202_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_176_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09106_ _04283_ _00715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_164_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06318_ _02173_ soc.spi_video_ram_1.write_fifo.fifo_mem\[18\]\[26\] _02119_ _02174_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xcaravel_hack_soc_206 wbs_dat_o[14] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
X_07298_ soc.spi_video_ram_1.write_fifo.fifo_mem\[18\]\[10\] soc.spi_video_ram_1.write_fifo.fifo_mem\[19\]\[10\]
+ _02893_ _02948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_87_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_191_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xcaravel_hack_soc_217 wbs_dat_o[25] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xcaravel_hack_soc_228 io_oeb[33] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
X_09037_ _04242_ _00687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_163_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06249_ _02127_ _00015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_102_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_46_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_213_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09939_ _04834_ _04838_ _04842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_24_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_245_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_234_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11901_ _00960_ clknet_leaf_44_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[3\]\[27\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_245_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_172_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_46_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11832_ _00891_ clknet_leaf_125_wb_clk_i soc.rom_encoder_0.input_buffer\[6\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1810 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1821 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_304_wb_clk_i clknet_5_1_0_wb_clk_i clknet_leaf_304_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_1832 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_226_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1843 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1854 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11763_ _00824_ clknet_leaf_68_wb_clk_i soc.spi_video_ram_1.state_sram_clk_counter\[6\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffnq_1
XFILLER_42_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1865 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_187_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_159_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10714_ soc.spi_video_ram_1.fifo_in_address\[8\] _05325_ _05338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_1887 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1898 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11694_ _00755_ clknet_leaf_304_wb_clk_i soc.spi_video_ram_1.fifo_in_data\[12\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_105_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_220_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_161_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10645_ soc.spi_video_ram_1.write_fifo.fifo_mem\[19\]\[21\] _04061_ _05277_ _05301_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_155_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_154_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10576_ soc.cpu.AReg.data\[0\] _01455_ _01572_ _01641_ _05261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_182_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12315_ _01343_ clknet_leaf_117_wb_clk_i soc.ram_encoder_0.data_out\[10\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_115_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_237_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12246_ _01274_ clknet_leaf_304_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[29\]\[28\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_218_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_159_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12177_ _01205_ clknet_leaf_85_wb_clk_i soc.boot_loading_offset\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_64_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_20_wb_clk_i clknet_5_2_0_wb_clk_i clknet_leaf_20_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_111_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_1_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_155_1398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_150_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11128_ _00194_ clknet_leaf_176_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[14\]\[8\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_228_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5170 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11059_ _00125_ clknet_leaf_293_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[0\]\[26\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_5181 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_224_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05620_ _01471_ _01528_ _01529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_92_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_240_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3790 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_166_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05551_ soc.spi_video_ram_1.buffer_index\[4\] _01460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_178_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_220_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08270_ soc.ram_encoder_0.output_buffer\[14\] _03814_ _03789_ soc.ram_encoder_0.request_data_out\[10\]
+ _03817_ _03825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_32_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05482_ _01393_ _01397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_149_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07221_ soc.spi_video_ram_1.write_fifo.fifo_mem\[24\]\[8\] soc.spi_video_ram_1.write_fifo.fifo_mem\[25\]\[8\]
+ soc.spi_video_ram_1.write_fifo.fifo_mem\[26\]\[8\] soc.spi_video_ram_1.write_fifo.fifo_mem\[27\]\[8\]
+ _02607_ _02578_ _02873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_203_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07152_ _02643_ _02806_ _02807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_140_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_173_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06103_ soc.video_generator_1.h_count\[1\] _01994_ _01995_ _01996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_145_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07083_ _02576_ _02740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_118_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_156_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_06034_ _01880_ _01888_ _01855_ _01876_ _01927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_161_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_216_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_232_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07985_ _03618_ _03620_ _03622_ _03624_ _02710_ _03625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_09724_ _04676_ _04678_ _04688_ _01381_ _00929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_80_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_210_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06936_ _02590_ _02597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_86_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_227_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_216_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09655_ _04636_ _00912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_28_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06867_ _01682_ _02534_ _02536_ _02537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_243_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08606_ _04007_ _00491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_83_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_05818_ _01563_ _01570_ _01718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_09586_ soc.rom_encoder_0.input_buffer\[3\] _04592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_27_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06798_ soc.rom_encoder_0.output_buffer\[19\] _02455_ _02474_ _02461_ _02475_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XTAP_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08537_ _02126_ soc.spi_video_ram_1.write_fifo.fifo_mem\[2\]\[3\] _03967_ _03971_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_05749_ _01595_ _01652_ _01653_ soc.cpu.PC.in\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_70_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_208_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_243_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_1488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_196_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08468_ _03933_ _03934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_51_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07419_ _03041_ _03064_ _03067_ _02570_ _03068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_221_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08399_ _03895_ _00396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_104_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_177_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10430_ _01615_ _01751_ _05157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_178_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_100_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10361_ _01834_ _05104_ _05120_ _01134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_30_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12100_ _01128_ net85 soc.cpu.ALU.x\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_139_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10292_ _05071_ _05077_ _05078_ _01106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_219_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_152_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_12031_ _01090_ clknet_leaf_72_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[5\]\[19\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_156_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_239_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3020 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3031 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_206_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3042 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3053 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xcaravel_hack_soc_93 io_oeb[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_74_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3064 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3075 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_233_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_185_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3086 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_222_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3097 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11815_ _00874_ clknet_leaf_48_wb_clk_i soc.spi_video_ram_1.write_fifo.write_pointer\[2\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_202_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_11746_ _00807_ clknet_leaf_70_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[4\]\[19\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_30_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1695 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_186_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11677_ _00738_ clknet_leaf_64_wb_clk_i soc.video_generator_1.v_count\[5\] vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_70_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10628_ _05292_ _01229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_200_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_155_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_239_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_196_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_182_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10559_ soc.boot_loading_offset\[2\] soc.boot_loading_offset\[1\] _05246_ _05250_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_143_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_155_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_185_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12229_ _01257_ clknet_leaf_36_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[29\]\[11\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_190_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_155_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_233_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_229_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_151_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_297_wb_clk_i clknet_5_4_0_wb_clk_i clknet_leaf_297_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_81_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07770_ soc.spi_video_ram_1.write_fifo.fifo_mem\[0\]\[15\] soc.spi_video_ram_1.write_fifo.fifo_mem\[1\]\[15\]
+ soc.spi_video_ram_1.write_fifo.fifo_mem\[2\]\[15\] soc.spi_video_ram_1.write_fifo.fifo_mem\[3\]\[15\]
+ _03139_ _02895_ _03415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_211_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_209_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_226_wb_clk_i clknet_5_21_0_wb_clk_i clknet_leaf_226_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_133_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_06721_ _02416_ _00198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_225_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09440_ soc.rom_encoder_0.request_address\[12\] _02520_ _04460_ soc.rom_encoder_0.output_buffer\[9\]
+ _04490_ _04491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_0_1713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06652_ _02151_ soc.spi_video_ram_1.write_fifo.fifo_mem\[12\]\[15\] _02368_ _02374_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_77_1439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05603_ _01473_ _01511_ _01512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_75_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09371_ soc.spi_video_ram_1.state_sram_clk_counter\[4\] _04439_ _04433_ _04442_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06583_ soc.spi_video_ram_1.write_fifo.fifo_mem\[13\]\[15\] _02248_ _02328_ _02334_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_80_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_209_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08322_ _02163_ soc.spi_video_ram_1.write_fifo.fifo_mem\[1\]\[21\] _03830_ _03854_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_05534_ _01405_ _01444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_221_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_178_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_240_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08253_ soc.ram_encoder_0.output_buffer\[11\] _03780_ _03811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_05465_ _01380_ _01381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_123_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_222_1753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07204_ soc.spi_video_ram_1.write_fifo.fifo_mem\[0\]\[7\] soc.spi_video_ram_1.write_fifo.fifo_mem\[1\]\[7\]
+ soc.spi_video_ram_1.write_fifo.fifo_mem\[2\]\[7\] soc.spi_video_ram_1.write_fifo.fifo_mem\[3\]\[7\]
+ _02680_ _02838_ _02857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_08184_ _02169_ soc.spi_video_ram_1.write_fifo.fifo_mem\[10\]\[24\] _03731_ _03758_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_118_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_146_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07135_ _02710_ _02781_ _02790_ _02791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_119_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_238_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07066_ _02697_ soc.spi_video_ram_1.write_fifo.fifo_mem\[31\]\[2\] _02725_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_133_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_245_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_06017_ _01885_ _01858_ _01868_ _01909_ _01910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_121_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_245_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_160_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5906 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_47_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_5917 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_88_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_1284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5928 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_87_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5939 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_1410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_74_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07968_ soc.spi_video_ram_1.write_fifo.fifo_mem\[28\]\[19\] soc.spi_video_ram_1.write_fifo.fifo_mem\[29\]\[19\]
+ soc.spi_video_ram_1.write_fifo.fifo_mem\[30\]\[19\] soc.spi_video_ram_1.write_fifo.fifo_mem\[31\]\[19\]
+ _02701_ _02737_ _03609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_114_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_1465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09707_ _04673_ _00927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06919_ _02571_ _02579_ _02580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_112_1544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07899_ _02645_ _03541_ _03542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_74_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09638_ _04627_ _00904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_112_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_215_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_204_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_186_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09569_ _04568_ _04577_ _04580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_167_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11600_ _00666_ clknet_leaf_194_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[21\]\[7\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_145_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_180_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_211_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_168_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_157_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11531_ _00597_ clknet_leaf_242_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[23\]\[25\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_54_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_1550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_184_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11462_ _00528_ clknet_leaf_309_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[15\]\[14\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_137_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_165_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10413_ _05148_ _01158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_109_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_183_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_164_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11393_ _00459_ clknet_leaf_259_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[2\]\[3\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_87_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_152_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_178_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_174_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10344_ soc.cpu.ALU.x\[6\] _05109_ _05112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_180_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_174_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_155_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10275_ soc.rom_loader.writing soc.rom_loader.was_loading _04611_ _05068_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_191_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12014_ _01073_ clknet_leaf_266_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[5\]\[2\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_61_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_215_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_238_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_207_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_189_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_47_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2160 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2171 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2182 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_203_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_241_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_187_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_163_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11729_ _00790_ clknet_leaf_254_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[4\]\[2\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_30_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_204_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_171_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_183_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_239_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_115_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_170_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_157_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08940_ _04191_ _00641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_142_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08871_ soc.spi_video_ram_1.write_fifo.fifo_mem\[25\]\[9\] _02409_ _04144_ _04154_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_170_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07822_ _02931_ soc.spi_video_ram_1.write_fifo.fifo_mem\[12\]\[23\] _03467_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_57_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07753_ _02752_ soc.spi_video_ram_1.write_fifo.fifo_mem\[28\]\[15\] _03397_ _02927_
+ _03398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_42_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06704_ soc.spi_video_ram_1.fifo_in_data\[7\] _02405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_07684_ soc.spi_video_ram_1.write_fifo.fifo_mem\[18\]\[24\] soc.spi_video_ram_1.write_fifo.fifo_mem\[19\]\[24\]
+ _02612_ _03330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_77_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_246_1539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09423_ soc.rom_encoder_0.request_address\[8\] _02520_ _04460_ soc.rom_encoder_0.output_buffer\[5\]
+ _04477_ _04478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_38_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06635_ _02134_ soc.spi_video_ram_1.write_fifo.fifo_mem\[12\]\[7\] _02357_ _02365_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_168_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_244_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_240_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09354_ _04428_ _04295_ _04429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_40_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06566_ soc.spi_video_ram_1.write_fifo.fifo_mem\[13\]\[7\] _02231_ _02317_ _02325_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_181_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08305_ _03845_ _00352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_107_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_05517_ _01430_ soc.spi_video_ram_1.current_state\[2\] _01431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_09285_ _02274_ soc.spi_video_ram_1.write_fifo.fifo_mem\[9\]\[28\] _04359_ _04391_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_139_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06497_ _02132_ soc.spi_video_ram_1.write_fifo.fifo_mem\[0\]\[6\] _02279_ _02286_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_166_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08236_ _02556_ _03797_ _03798_ _00330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_53_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_165_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08167_ _03749_ _00310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_119_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_146_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_175_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_1245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07118_ _01534_ _02676_ _02735_ _02774_ _00236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_179_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08098_ _03708_ _00282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_175_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_162_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07049_ _02693_ _02699_ _02702_ _02705_ _02707_ _02708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XTAP_6415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_6437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_148_wb_clk_i clknet_5_28_0_wb_clk_i clknet_leaf_148_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_134_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_6448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5703 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10060_ soc.ram_encoder_0.initializing_step\[3\] _04916_ _04684_ _04917_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_6459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5714 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_138_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5725 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5736 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5747 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5758 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_130_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5769 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_153_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_188_1718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_169_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_244_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10962_ _00028_ clknet_leaf_79_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[18\]\[16\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_44_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_243_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10893_ soc.spi_video_ram_1.write_fifo.fifo_mem\[8\]\[3\] soc.spi_video_ram_1.fifo_in_data\[3\]
+ _05431_ _05435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_232_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_145_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_169_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_145_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11514_ _00580_ clknet_leaf_208_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[23\]\[8\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_7_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12494_ net57 net54 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_221_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11445_ _00511_ clknet_leaf_294_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[30\]\[26\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_32_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11376_ _00442_ clknet_leaf_311_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[28\]\[15\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_113_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_153_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10327_ soc.rom_loader.wait_fall_clk _05100_ _05101_ _01118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_152_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_158_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_106_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_234_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10258_ _03453_ _05044_ _05057_ _01094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_26_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_152_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_45_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_152_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_239_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10189_ soc.hack_clock_0.counter\[1\] soc.hack_clock_0.counter\[0\] _05018_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_26_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_212_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_152_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_187_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_234_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06420_ soc.spi_video_ram_1.fifo_in_data\[9\] _02235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_222_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_245_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_98_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_50_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_163_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06351_ _02140_ soc.spi_video_ram_1.write_fifo.fifo_mem\[17\]\[10\] _02193_ _02194_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_30_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_148_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09070_ _02227_ soc.spi_video_ram_1.write_fifo.fifo_mem\[20\]\[5\] _04259_ _04265_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_136_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06282_ _02149_ soc.spi_video_ram_1.write_fifo.fifo_mem\[18\]\[14\] _02141_ _02150_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_124_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08021_ soc.spi_video_ram_1.write_fifo.fifo_mem\[4\]\[16\] soc.spi_video_ram_1.write_fifo.fifo_mem\[5\]\[16\]
+ soc.spi_video_ram_1.write_fifo.fifo_mem\[6\]\[16\] soc.spi_video_ram_1.write_fifo.fifo_mem\[7\]\[16\]
+ _02701_ _03041_ _03659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_11_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_198_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_200_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_157_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_171_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09972_ soc.ram_encoder_0.input_buffer\[8\] _04865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_118_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_241_wb_clk_i clknet_5_16_0_wb_clk_i clknet_leaf_241_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_08923_ _04182_ _00633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_44_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_130_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08854_ _04145_ _00601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_170_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_1279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_57_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07805_ soc.spi_video_ram_1.write_fifo.fifo_mem\[7\]\[23\] _03450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_3608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08785_ _04106_ _00571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_05997_ _01876_ _01889_ _01890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_73_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_226_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_211_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2907 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07736_ _03047_ soc.spi_video_ram_1.write_fifo.fifo_mem\[17\]\[15\] _03381_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_77_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2918 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2929 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_246_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_164_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07667_ _02644_ _03312_ _03313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_246_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_225_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_214_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09406_ soc.rom_encoder_0.output_buffer\[2\] _04460_ _04464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_06618_ _02116_ _02214_ _02313_ _02355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_164_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_241_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_198_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07598_ soc.spi_video_ram_1.write_fifo.fifo_mem\[24\]\[25\] soc.spi_video_ram_1.write_fifo.fifo_mem\[25\]\[25\]
+ soc.spi_video_ram_1.write_fifo.fifo_mem\[26\]\[25\] soc.spi_video_ram_1.write_fifo.fifo_mem\[27\]\[25\]
+ _02907_ _02908_ _03245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_142_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09337_ _04419_ _00810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06549_ _02311_ _02314_ _02315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_55_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_224_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09268_ _04382_ _00778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_127_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_194_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08219_ _02556_ _03784_ _03785_ _00326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_177_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09199_ soc.spi_video_ram_1.fifo_in_data\[4\] _04341_ _04345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_5_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11230_ _00296_ clknet_leaf_205_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[10\]\[1\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_88_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_162_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_155_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_150_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11161_ _00227_ clknet_leaf_105_wb_clk_i soc.rom_encoder_0.output_buffer\[2\] vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_6201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_235_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_6212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10112_ _04855_ _04947_ _04948_ _04959_ _04960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_6234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_175_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_6245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11092_ _00158_ clknet_leaf_224_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[12\]\[1\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_110_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_88_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_216_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10043_ _04907_ _01029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_6289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_1357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4810 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_130_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4821 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_5577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4832 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_5588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4843 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4854 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4865 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4876 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_29_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4887 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_1_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4898 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_99_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11994_ _01053_ clknet_leaf_118_wb_clk_i soc.ram_data_out\[15\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_216_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_72_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10945_ _05461_ _01377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_43_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_45_wb_clk_i clknet_5_6_0_wb_clk_i clknet_leaf_45_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_204_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_177_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_147_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10876_ soc.ram_encoder_0.data_out\[12\] _05425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_143_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_242_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_227_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_231_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_188_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_164_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_77_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_200_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_145_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_184_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_199_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_4 _05266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_201_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11428_ _00494_ clknet_leaf_255_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[30\]\[9\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_126_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_158_1352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_153_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11359_ _00425_ clknet_leaf_297_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[27\]\[27\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_98_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_193_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_154_1249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_05920_ _01786_ _01813_ _01814_ _01815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_67_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_05851_ _01682_ _01740_ _01743_ _01750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_13_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_208_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_187_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08570_ _02159_ soc.spi_video_ram_1.write_fifo.fifo_mem\[2\]\[19\] _03978_ _03988_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_05782_ _01557_ _01683_ _01684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_235_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07521_ soc.spi_video_ram_1.write_fifo.fifo_mem\[15\]\[26\] _03169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_207_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07452_ _02567_ _03093_ _03100_ _03101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_223_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_161_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_228_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06403_ soc.spi_video_ram_1.write_fifo.fifo_mem\[16\]\[3\] _02223_ _02217_ _02224_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_182_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_194_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07383_ _02719_ _03026_ _03031_ _03032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_91_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09122_ _01414_ _04292_ _01379_ _04293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_06334_ _02124_ soc.spi_video_ram_1.write_fifo.fifo_mem\[17\]\[2\] _02182_ _02185_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_206_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_241_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_148_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09053_ _01380_ _04254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_11_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_148_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06265_ soc.spi_video_ram_1.fifo_in_data\[9\] _02138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_136_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08004_ soc.spi_video_ram_1.write_fifo.fifo_mem\[4\]\[17\] soc.spi_video_ram_1.write_fifo.fifo_mem\[5\]\[17\]
+ soc.spi_video_ram_1.write_fifo.fifo_mem\[6\]\[17\] soc.spi_video_ram_1.write_fifo.fifo_mem\[7\]\[17\]
+ _02717_ _02682_ _03643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_159_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_219_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_191_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06196_ _01520_ _01523_ _02083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_89_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_176_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_219_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09955_ net3 _04849_ _04601_ _04854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_106_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_217_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08906_ soc.spi_video_ram_1.write_fifo.fifo_mem\[25\]\[26\] _03927_ _04143_ _04172_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_4106 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09886_ _04738_ _04800_ net62 _04801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4117 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_4128 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_170_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_4139 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08837_ _03482_ _04124_ _04135_ _00594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_3405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_246_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2704 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08768_ soc.spi_video_ram_1.write_fifo.fifo_mem\[24\]\[20\] _02343_ _04075_ _04098_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_2715 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2726 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_245_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_26_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2737 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_148_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_246_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07719_ _02679_ _03364_ _03365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_57_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2748 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2759 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08699_ soc.spi_video_ram_1.write_fifo.fifo_mem\[15\]\[19\] _02341_ _04043_ _04059_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_41_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_198_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10730_ soc.spi_video_ram_1.write_fifo.fifo_mem\[31\]\[2\] soc.spi_video_ram_1.fifo_in_data\[2\]
+ _05344_ _05347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_199_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_213_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10661_ _03931_ _02179_ _05309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_161_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_210_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10592_ _05270_ _05268_ _05271_ _01214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_107_1284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12331_ _01359_ clknet_leaf_13_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[8\]\[10\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_215_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_166_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_163_wb_clk_i clknet_5_27_0_wb_clk_i clknet_leaf_163_wb_clk_i vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_12262_ _01290_ clknet_leaf_311_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[31\]\[15\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_182_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11213_ _00279_ clknet_leaf_238_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[11\]\[23\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_135_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12193_ _01221_ clknet_leaf_139_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[19\]\[4\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_107_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput52 net52 io_oeb[18] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_194_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11144_ _00210_ clknet_leaf_306_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[14\]\[24\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_6020 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput63 net63 io_out[15] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_6031 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput74 net74 io_out[27] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_96_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_6042 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6053 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6064 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_150_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11075_ _00141_ clknet_leaf_16_wb_clk_i soc.spi_video_ram_1.write_fifo.fifo_mem\[13\]\[13\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_6075 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_163_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_6086 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_6097 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_5363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10026_ _04898_ _01021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_76_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_5374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_188_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_5385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_4651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_5396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_4662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_4673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_4695 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3950 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_236_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3961 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_217_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3972 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3983 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11977_ _01036_ clknet_leaf_153_wb_clk_i soc.ram_encoder_0.request_address\[14\]
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_3994 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_225_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_205_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10928_ soc.spi_video_ram_1.write_fifo.fifo_mem\[8\]\[20\] soc.spi_video_ram_1.fifo_in_address\[4\]
+ _05430_ _05453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_176_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_147_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_189_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10859_ _01652_ _05222_ _05412_ _05416_ _01336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_125_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_34_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_173_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_201_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_158_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_173_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06050_ _01868_ _01928_ _01929_ _01935_ _01943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_133_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_207_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_236_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06952_ _02612_ _02613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
X_09740_ _04699_ _00934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_100_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
.ends

